// This is the unpowered netlist.
module wrapped_as2650 (wb_clk_i,
    io_in,
    io_oeb,
    io_out);
 input wb_clk_i;
 input [37:0] io_in;
 output [37:0] io_oeb;
 output [37:0] io_out;

 wire net85;
 wire net90;
 wire net55;
 wire net56;
 wire net57;
 wire net58;
 wire net59;
 wire net60;
 wire net86;
 wire net61;
 wire net62;
 wire net63;
 wire net64;
 wire net65;
 wire net66;
 wire net67;
 wire net68;
 wire net69;
 wire net70;
 wire net87;
 wire net71;
 wire net72;
 wire net73;
 wire net91;
 wire net92;
 wire net93;
 wire net94;
 wire net95;
 wire net88;
 wire net89;
 wire net74;
 wire net79;
 wire net75;
 wire net76;
 wire net80;
 wire net81;
 wire net82;
 wire net83;
 wire net84;
 wire net77;
 wire net78;
 wire _0000_;
 wire _0001_;
 wire _0002_;
 wire _0003_;
 wire _0004_;
 wire _0005_;
 wire _0006_;
 wire _0007_;
 wire _0008_;
 wire _0009_;
 wire _0010_;
 wire _0011_;
 wire _0012_;
 wire _0013_;
 wire _0014_;
 wire _0015_;
 wire _0016_;
 wire _0017_;
 wire _0018_;
 wire _0019_;
 wire _0020_;
 wire _0021_;
 wire _0022_;
 wire _0023_;
 wire _0024_;
 wire _0025_;
 wire _0026_;
 wire _0027_;
 wire _0028_;
 wire _0029_;
 wire _0030_;
 wire _0031_;
 wire _0032_;
 wire _0033_;
 wire _0034_;
 wire _0035_;
 wire _0036_;
 wire _0037_;
 wire _0038_;
 wire _0039_;
 wire _0040_;
 wire _0041_;
 wire _0042_;
 wire _0043_;
 wire _0044_;
 wire _0045_;
 wire _0046_;
 wire _0047_;
 wire _0048_;
 wire _0049_;
 wire _0050_;
 wire _0051_;
 wire _0052_;
 wire _0053_;
 wire _0054_;
 wire _0055_;
 wire _0056_;
 wire _0057_;
 wire _0058_;
 wire _0059_;
 wire _0060_;
 wire _0061_;
 wire _0062_;
 wire _0063_;
 wire _0064_;
 wire _0065_;
 wire _0066_;
 wire _0067_;
 wire _0068_;
 wire _0069_;
 wire _0070_;
 wire _0071_;
 wire _0072_;
 wire _0073_;
 wire _0074_;
 wire _0075_;
 wire _0076_;
 wire _0077_;
 wire _0078_;
 wire _0079_;
 wire _0080_;
 wire _0081_;
 wire _0082_;
 wire _0083_;
 wire _0084_;
 wire _0085_;
 wire _0086_;
 wire _0087_;
 wire _0088_;
 wire _0089_;
 wire _0090_;
 wire _0091_;
 wire _0092_;
 wire _0093_;
 wire _0094_;
 wire _0095_;
 wire _0096_;
 wire _0097_;
 wire _0098_;
 wire _0099_;
 wire _0100_;
 wire _0101_;
 wire _0102_;
 wire _0103_;
 wire _0104_;
 wire _0105_;
 wire _0106_;
 wire _0107_;
 wire _0108_;
 wire _0109_;
 wire _0110_;
 wire _0111_;
 wire _0112_;
 wire _0113_;
 wire _0114_;
 wire _0115_;
 wire _0116_;
 wire _0117_;
 wire _0118_;
 wire _0119_;
 wire _0120_;
 wire _0121_;
 wire _0122_;
 wire _0123_;
 wire _0124_;
 wire _0125_;
 wire _0126_;
 wire _0127_;
 wire _0128_;
 wire _0129_;
 wire _0130_;
 wire _0131_;
 wire _0132_;
 wire _0133_;
 wire _0134_;
 wire _0135_;
 wire _0136_;
 wire _0137_;
 wire _0138_;
 wire _0139_;
 wire _0140_;
 wire _0141_;
 wire _0142_;
 wire _0143_;
 wire _0144_;
 wire _0145_;
 wire _0146_;
 wire _0147_;
 wire _0148_;
 wire _0149_;
 wire _0150_;
 wire _0151_;
 wire _0152_;
 wire _0153_;
 wire _0154_;
 wire _0155_;
 wire _0156_;
 wire _0157_;
 wire _0158_;
 wire _0159_;
 wire _0160_;
 wire _0161_;
 wire _0162_;
 wire _0163_;
 wire _0164_;
 wire _0165_;
 wire _0166_;
 wire _0167_;
 wire _0168_;
 wire _0169_;
 wire _0170_;
 wire _0171_;
 wire _0172_;
 wire _0173_;
 wire _0174_;
 wire _0175_;
 wire _0176_;
 wire _0177_;
 wire _0178_;
 wire _0179_;
 wire _0180_;
 wire _0181_;
 wire _0182_;
 wire _0183_;
 wire _0184_;
 wire _0185_;
 wire _0186_;
 wire _0187_;
 wire _0188_;
 wire _0189_;
 wire _0190_;
 wire _0191_;
 wire _0192_;
 wire _0193_;
 wire _0194_;
 wire _0195_;
 wire _0196_;
 wire _0197_;
 wire _0198_;
 wire _0199_;
 wire _0200_;
 wire _0201_;
 wire _0202_;
 wire _0203_;
 wire _0204_;
 wire _0205_;
 wire _0206_;
 wire _0207_;
 wire _0208_;
 wire _0209_;
 wire _0210_;
 wire _0211_;
 wire _0212_;
 wire _0213_;
 wire _0214_;
 wire _0215_;
 wire _0216_;
 wire _0217_;
 wire _0218_;
 wire _0219_;
 wire _0220_;
 wire _0221_;
 wire _0222_;
 wire _0223_;
 wire _0224_;
 wire _0225_;
 wire _0226_;
 wire _0227_;
 wire _0228_;
 wire _0229_;
 wire _0230_;
 wire _0231_;
 wire _0232_;
 wire _0233_;
 wire _0234_;
 wire _0235_;
 wire _0236_;
 wire _0237_;
 wire _0238_;
 wire _0239_;
 wire _0240_;
 wire _0241_;
 wire _0242_;
 wire _0243_;
 wire _0244_;
 wire _0245_;
 wire _0246_;
 wire _0247_;
 wire _0248_;
 wire _0249_;
 wire _0250_;
 wire _0251_;
 wire _0252_;
 wire _0253_;
 wire _0254_;
 wire _0255_;
 wire _0256_;
 wire _0257_;
 wire _0258_;
 wire _0259_;
 wire _0260_;
 wire _0261_;
 wire _0262_;
 wire _0263_;
 wire _0264_;
 wire _0265_;
 wire _0266_;
 wire _0267_;
 wire _0268_;
 wire _0269_;
 wire _0270_;
 wire _0271_;
 wire _0272_;
 wire _0273_;
 wire _0274_;
 wire _0275_;
 wire _0276_;
 wire _0277_;
 wire _0278_;
 wire _0279_;
 wire _0280_;
 wire _0281_;
 wire _0282_;
 wire _0283_;
 wire _0284_;
 wire _0285_;
 wire _0286_;
 wire _0287_;
 wire _0288_;
 wire _0289_;
 wire _0290_;
 wire _0291_;
 wire _0292_;
 wire _0293_;
 wire _0294_;
 wire _0295_;
 wire _0296_;
 wire _0297_;
 wire _0298_;
 wire _0299_;
 wire _0300_;
 wire _0301_;
 wire _0302_;
 wire _0303_;
 wire _0304_;
 wire _0305_;
 wire _0306_;
 wire _0307_;
 wire _0308_;
 wire _0309_;
 wire _0310_;
 wire _0311_;
 wire _0312_;
 wire _0313_;
 wire _0314_;
 wire _0315_;
 wire _0316_;
 wire _0317_;
 wire _0318_;
 wire _0319_;
 wire _0320_;
 wire _0321_;
 wire _0322_;
 wire _0323_;
 wire _0324_;
 wire _0325_;
 wire _0326_;
 wire _0327_;
 wire _0328_;
 wire _0329_;
 wire _0330_;
 wire _0331_;
 wire _0332_;
 wire _0333_;
 wire _0334_;
 wire _0335_;
 wire _0336_;
 wire _0337_;
 wire _0338_;
 wire _0339_;
 wire _0340_;
 wire _0341_;
 wire _0342_;
 wire _0343_;
 wire _0344_;
 wire _0345_;
 wire _0346_;
 wire _0347_;
 wire _0348_;
 wire _0349_;
 wire _0350_;
 wire _0351_;
 wire _0352_;
 wire _0353_;
 wire _0354_;
 wire _0355_;
 wire _0356_;
 wire _0357_;
 wire _0358_;
 wire _0359_;
 wire _0360_;
 wire _0361_;
 wire _0362_;
 wire _0363_;
 wire _0364_;
 wire _0365_;
 wire _0366_;
 wire _0367_;
 wire _0368_;
 wire _0369_;
 wire _0370_;
 wire _0371_;
 wire _0372_;
 wire _0373_;
 wire _0374_;
 wire _0375_;
 wire _0376_;
 wire _0377_;
 wire _0378_;
 wire _0379_;
 wire _0380_;
 wire _0381_;
 wire _0382_;
 wire _0383_;
 wire _0384_;
 wire _0385_;
 wire _0386_;
 wire _0387_;
 wire _0388_;
 wire _0389_;
 wire _0390_;
 wire _0391_;
 wire _0392_;
 wire _0393_;
 wire _0394_;
 wire _0395_;
 wire _0396_;
 wire _0397_;
 wire _0398_;
 wire _0399_;
 wire _0400_;
 wire _0401_;
 wire _0402_;
 wire _0403_;
 wire _0404_;
 wire _0405_;
 wire _0406_;
 wire _0407_;
 wire _0408_;
 wire _0409_;
 wire _0410_;
 wire _0411_;
 wire _0412_;
 wire _0413_;
 wire _0414_;
 wire _0415_;
 wire _0416_;
 wire _0417_;
 wire _0418_;
 wire _0419_;
 wire _0420_;
 wire _0421_;
 wire _0422_;
 wire _0423_;
 wire _0424_;
 wire _0425_;
 wire _0426_;
 wire _0427_;
 wire _0428_;
 wire _0429_;
 wire _0430_;
 wire _0431_;
 wire _0432_;
 wire _0433_;
 wire _0434_;
 wire _0435_;
 wire _0436_;
 wire _0437_;
 wire _0438_;
 wire _0439_;
 wire _0440_;
 wire _0441_;
 wire _0442_;
 wire _0443_;
 wire _0444_;
 wire _0445_;
 wire _0446_;
 wire _0447_;
 wire _0448_;
 wire _0449_;
 wire _0450_;
 wire _0451_;
 wire _0452_;
 wire _0453_;
 wire _0454_;
 wire _0455_;
 wire _0456_;
 wire _0457_;
 wire _0458_;
 wire _0459_;
 wire _0460_;
 wire _0461_;
 wire _0462_;
 wire _0463_;
 wire _0464_;
 wire _0465_;
 wire _0466_;
 wire _0467_;
 wire _0468_;
 wire _0469_;
 wire _0470_;
 wire _0471_;
 wire _0472_;
 wire _0473_;
 wire _0474_;
 wire _0475_;
 wire _0476_;
 wire _0477_;
 wire _0478_;
 wire _0479_;
 wire _0480_;
 wire _0481_;
 wire _0482_;
 wire _0483_;
 wire _0484_;
 wire _0485_;
 wire _0486_;
 wire _0487_;
 wire _0488_;
 wire _0489_;
 wire _0490_;
 wire _0491_;
 wire _0492_;
 wire _0493_;
 wire _0494_;
 wire _0495_;
 wire _0496_;
 wire _0497_;
 wire _0498_;
 wire _0499_;
 wire _0500_;
 wire _0501_;
 wire _0502_;
 wire _0503_;
 wire _0504_;
 wire _0505_;
 wire _0506_;
 wire _0507_;
 wire _0508_;
 wire _0509_;
 wire _0510_;
 wire _0511_;
 wire _0512_;
 wire _0513_;
 wire _0514_;
 wire _0515_;
 wire _0516_;
 wire _0517_;
 wire _0518_;
 wire _0519_;
 wire _0520_;
 wire _0521_;
 wire _0522_;
 wire _0523_;
 wire _0524_;
 wire _0525_;
 wire _0526_;
 wire _0527_;
 wire _0528_;
 wire _0529_;
 wire _0530_;
 wire _0531_;
 wire _0532_;
 wire _0533_;
 wire _0534_;
 wire _0535_;
 wire _0536_;
 wire _0537_;
 wire _0538_;
 wire _0539_;
 wire _0540_;
 wire _0541_;
 wire _0542_;
 wire _0543_;
 wire _0544_;
 wire _0545_;
 wire _0546_;
 wire _0547_;
 wire _0548_;
 wire _0549_;
 wire _0550_;
 wire _0551_;
 wire _0552_;
 wire _0553_;
 wire _0554_;
 wire _0555_;
 wire _0556_;
 wire _0557_;
 wire _0558_;
 wire _0559_;
 wire _0560_;
 wire _0561_;
 wire _0562_;
 wire _0563_;
 wire _0564_;
 wire _0565_;
 wire _0566_;
 wire _0567_;
 wire _0568_;
 wire _0569_;
 wire _0570_;
 wire _0571_;
 wire _0572_;
 wire _0573_;
 wire _0574_;
 wire _0575_;
 wire _0576_;
 wire _0577_;
 wire _0578_;
 wire _0579_;
 wire _0580_;
 wire _0581_;
 wire _0582_;
 wire _0583_;
 wire _0584_;
 wire _0585_;
 wire _0586_;
 wire _0587_;
 wire _0588_;
 wire _0589_;
 wire _0590_;
 wire _0591_;
 wire _0592_;
 wire _0593_;
 wire _0594_;
 wire _0595_;
 wire _0596_;
 wire _0597_;
 wire _0598_;
 wire _0599_;
 wire _0600_;
 wire _0601_;
 wire _0602_;
 wire _0603_;
 wire _0604_;
 wire _0605_;
 wire _0606_;
 wire _0607_;
 wire _0608_;
 wire _0609_;
 wire _0610_;
 wire _0611_;
 wire _0612_;
 wire _0613_;
 wire _0614_;
 wire _0615_;
 wire _0616_;
 wire _0617_;
 wire _0618_;
 wire _0619_;
 wire _0620_;
 wire _0621_;
 wire _0622_;
 wire _0623_;
 wire _0624_;
 wire _0625_;
 wire _0626_;
 wire _0627_;
 wire _0628_;
 wire _0629_;
 wire _0630_;
 wire _0631_;
 wire _0632_;
 wire _0633_;
 wire _0634_;
 wire _0635_;
 wire _0636_;
 wire _0637_;
 wire _0638_;
 wire _0639_;
 wire _0640_;
 wire _0641_;
 wire _0642_;
 wire _0643_;
 wire _0644_;
 wire _0645_;
 wire _0646_;
 wire _0647_;
 wire _0648_;
 wire _0649_;
 wire _0650_;
 wire _0651_;
 wire _0652_;
 wire _0653_;
 wire _0654_;
 wire _0655_;
 wire _0656_;
 wire _0657_;
 wire _0658_;
 wire _0659_;
 wire _0660_;
 wire _0661_;
 wire _0662_;
 wire _0663_;
 wire _0664_;
 wire _0665_;
 wire _0666_;
 wire _0667_;
 wire _0668_;
 wire _0669_;
 wire _0670_;
 wire _0671_;
 wire _0672_;
 wire _0673_;
 wire _0674_;
 wire _0675_;
 wire _0676_;
 wire _0677_;
 wire _0678_;
 wire _0679_;
 wire _0680_;
 wire _0681_;
 wire _0682_;
 wire _0683_;
 wire _0684_;
 wire _0685_;
 wire _0686_;
 wire _0687_;
 wire _0688_;
 wire _0689_;
 wire _0690_;
 wire _0691_;
 wire _0692_;
 wire _0693_;
 wire _0694_;
 wire _0695_;
 wire _0696_;
 wire _0697_;
 wire _0698_;
 wire _0699_;
 wire _0700_;
 wire _0701_;
 wire _0702_;
 wire _0703_;
 wire _0704_;
 wire _0705_;
 wire _0706_;
 wire _0707_;
 wire _0708_;
 wire _0709_;
 wire _0710_;
 wire _0711_;
 wire _0712_;
 wire _0713_;
 wire _0714_;
 wire _0715_;
 wire _0716_;
 wire _0717_;
 wire _0718_;
 wire _0719_;
 wire _0720_;
 wire _0721_;
 wire _0722_;
 wire _0723_;
 wire _0724_;
 wire _0725_;
 wire _0726_;
 wire _0727_;
 wire _0728_;
 wire _0729_;
 wire _0730_;
 wire _0731_;
 wire _0732_;
 wire _0733_;
 wire _0734_;
 wire _0735_;
 wire _0736_;
 wire _0737_;
 wire _0738_;
 wire _0739_;
 wire _0740_;
 wire _0741_;
 wire _0742_;
 wire _0743_;
 wire _0744_;
 wire _0745_;
 wire _0746_;
 wire _0747_;
 wire _0748_;
 wire _0749_;
 wire _0750_;
 wire _0751_;
 wire _0752_;
 wire _0753_;
 wire _0754_;
 wire _0755_;
 wire _0756_;
 wire _0757_;
 wire _0758_;
 wire _0759_;
 wire _0760_;
 wire _0761_;
 wire _0762_;
 wire _0763_;
 wire _0764_;
 wire _0765_;
 wire _0766_;
 wire _0767_;
 wire _0768_;
 wire _0769_;
 wire _0770_;
 wire _0771_;
 wire _0772_;
 wire _0773_;
 wire _0774_;
 wire _0775_;
 wire _0776_;
 wire _0777_;
 wire _0778_;
 wire _0779_;
 wire _0780_;
 wire _0781_;
 wire _0782_;
 wire _0783_;
 wire _0784_;
 wire _0785_;
 wire _0786_;
 wire _0787_;
 wire _0788_;
 wire _0789_;
 wire _0790_;
 wire _0791_;
 wire _0792_;
 wire _0793_;
 wire _0794_;
 wire _0795_;
 wire _0796_;
 wire _0797_;
 wire _0798_;
 wire _0799_;
 wire _0800_;
 wire _0801_;
 wire _0802_;
 wire _0803_;
 wire _0804_;
 wire _0805_;
 wire _0806_;
 wire _0807_;
 wire _0808_;
 wire _0809_;
 wire _0810_;
 wire _0811_;
 wire _0812_;
 wire _0813_;
 wire _0814_;
 wire _0815_;
 wire _0816_;
 wire _0817_;
 wire _0818_;
 wire _0819_;
 wire _0820_;
 wire _0821_;
 wire _0822_;
 wire _0823_;
 wire _0824_;
 wire _0825_;
 wire _0826_;
 wire _0827_;
 wire _0828_;
 wire _0829_;
 wire _0830_;
 wire _0831_;
 wire _0832_;
 wire _0833_;
 wire _0834_;
 wire _0835_;
 wire _0836_;
 wire _0837_;
 wire _0838_;
 wire _0839_;
 wire _0840_;
 wire _0841_;
 wire _0842_;
 wire _0843_;
 wire _0844_;
 wire _0845_;
 wire _0846_;
 wire _0847_;
 wire _0848_;
 wire _0849_;
 wire _0850_;
 wire _0851_;
 wire _0852_;
 wire _0853_;
 wire _0854_;
 wire _0855_;
 wire _0856_;
 wire _0857_;
 wire _0858_;
 wire _0859_;
 wire _0860_;
 wire _0861_;
 wire _0862_;
 wire _0863_;
 wire _0864_;
 wire _0865_;
 wire _0866_;
 wire _0867_;
 wire _0868_;
 wire _0869_;
 wire _0870_;
 wire _0871_;
 wire _0872_;
 wire _0873_;
 wire _0874_;
 wire _0875_;
 wire _0876_;
 wire _0877_;
 wire _0878_;
 wire _0879_;
 wire _0880_;
 wire _0881_;
 wire _0882_;
 wire _0883_;
 wire _0884_;
 wire _0885_;
 wire _0886_;
 wire _0887_;
 wire _0888_;
 wire _0889_;
 wire _0890_;
 wire _0891_;
 wire _0892_;
 wire _0893_;
 wire _0894_;
 wire _0895_;
 wire _0896_;
 wire _0897_;
 wire _0898_;
 wire _0899_;
 wire _0900_;
 wire _0901_;
 wire _0902_;
 wire _0903_;
 wire _0904_;
 wire _0905_;
 wire _0906_;
 wire _0907_;
 wire _0908_;
 wire _0909_;
 wire _0910_;
 wire _0911_;
 wire _0912_;
 wire _0913_;
 wire _0914_;
 wire _0915_;
 wire _0916_;
 wire _0917_;
 wire _0918_;
 wire _0919_;
 wire _0920_;
 wire _0921_;
 wire _0922_;
 wire _0923_;
 wire _0924_;
 wire _0925_;
 wire _0926_;
 wire _0927_;
 wire _0928_;
 wire _0929_;
 wire _0930_;
 wire _0931_;
 wire _0932_;
 wire _0933_;
 wire _0934_;
 wire _0935_;
 wire _0936_;
 wire _0937_;
 wire _0938_;
 wire _0939_;
 wire _0940_;
 wire _0941_;
 wire _0942_;
 wire _0943_;
 wire _0944_;
 wire _0945_;
 wire _0946_;
 wire _0947_;
 wire _0948_;
 wire _0949_;
 wire _0950_;
 wire _0951_;
 wire _0952_;
 wire _0953_;
 wire _0954_;
 wire _0955_;
 wire _0956_;
 wire _0957_;
 wire _0958_;
 wire _0959_;
 wire _0960_;
 wire _0961_;
 wire _0962_;
 wire _0963_;
 wire _0964_;
 wire _0965_;
 wire _0966_;
 wire _0967_;
 wire _0968_;
 wire _0969_;
 wire _0970_;
 wire _0971_;
 wire _0972_;
 wire _0973_;
 wire _0974_;
 wire _0975_;
 wire _0976_;
 wire _0977_;
 wire _0978_;
 wire _0979_;
 wire _0980_;
 wire _0981_;
 wire _0982_;
 wire _0983_;
 wire _0984_;
 wire _0985_;
 wire _0986_;
 wire _0987_;
 wire _0988_;
 wire _0989_;
 wire _0990_;
 wire _0991_;
 wire _0992_;
 wire _0993_;
 wire _0994_;
 wire _0995_;
 wire _0996_;
 wire _0997_;
 wire _0998_;
 wire _0999_;
 wire _1000_;
 wire _1001_;
 wire _1002_;
 wire _1003_;
 wire _1004_;
 wire _1005_;
 wire _1006_;
 wire _1007_;
 wire _1008_;
 wire _1009_;
 wire _1010_;
 wire _1011_;
 wire _1012_;
 wire _1013_;
 wire _1014_;
 wire _1015_;
 wire _1016_;
 wire _1017_;
 wire _1018_;
 wire _1019_;
 wire _1020_;
 wire _1021_;
 wire _1022_;
 wire _1023_;
 wire _1024_;
 wire _1025_;
 wire _1026_;
 wire _1027_;
 wire _1028_;
 wire _1029_;
 wire _1030_;
 wire _1031_;
 wire _1032_;
 wire _1033_;
 wire _1034_;
 wire _1035_;
 wire _1036_;
 wire _1037_;
 wire _1038_;
 wire _1039_;
 wire _1040_;
 wire _1041_;
 wire _1042_;
 wire _1043_;
 wire _1044_;
 wire _1045_;
 wire _1046_;
 wire _1047_;
 wire _1048_;
 wire _1049_;
 wire _1050_;
 wire _1051_;
 wire _1052_;
 wire _1053_;
 wire _1054_;
 wire _1055_;
 wire _1056_;
 wire _1057_;
 wire _1058_;
 wire _1059_;
 wire _1060_;
 wire _1061_;
 wire _1062_;
 wire _1063_;
 wire _1064_;
 wire _1065_;
 wire _1066_;
 wire _1067_;
 wire _1068_;
 wire _1069_;
 wire _1070_;
 wire _1071_;
 wire _1072_;
 wire _1073_;
 wire _1074_;
 wire _1075_;
 wire _1076_;
 wire _1077_;
 wire _1078_;
 wire _1079_;
 wire _1080_;
 wire _1081_;
 wire _1082_;
 wire _1083_;
 wire _1084_;
 wire _1085_;
 wire _1086_;
 wire _1087_;
 wire _1088_;
 wire _1089_;
 wire _1090_;
 wire _1091_;
 wire _1092_;
 wire _1093_;
 wire _1094_;
 wire _1095_;
 wire _1096_;
 wire _1097_;
 wire _1098_;
 wire _1099_;
 wire _1100_;
 wire _1101_;
 wire _1102_;
 wire _1103_;
 wire _1104_;
 wire _1105_;
 wire _1106_;
 wire _1107_;
 wire _1108_;
 wire _1109_;
 wire _1110_;
 wire _1111_;
 wire _1112_;
 wire _1113_;
 wire _1114_;
 wire _1115_;
 wire _1116_;
 wire _1117_;
 wire _1118_;
 wire _1119_;
 wire _1120_;
 wire _1121_;
 wire _1122_;
 wire _1123_;
 wire _1124_;
 wire _1125_;
 wire _1126_;
 wire _1127_;
 wire _1128_;
 wire _1129_;
 wire _1130_;
 wire _1131_;
 wire _1132_;
 wire _1133_;
 wire _1134_;
 wire _1135_;
 wire _1136_;
 wire _1137_;
 wire _1138_;
 wire _1139_;
 wire _1140_;
 wire _1141_;
 wire _1142_;
 wire _1143_;
 wire _1144_;
 wire _1145_;
 wire _1146_;
 wire _1147_;
 wire _1148_;
 wire _1149_;
 wire _1150_;
 wire _1151_;
 wire _1152_;
 wire _1153_;
 wire _1154_;
 wire _1155_;
 wire _1156_;
 wire _1157_;
 wire _1158_;
 wire _1159_;
 wire _1160_;
 wire _1161_;
 wire _1162_;
 wire _1163_;
 wire _1164_;
 wire _1165_;
 wire _1166_;
 wire _1167_;
 wire _1168_;
 wire _1169_;
 wire _1170_;
 wire _1171_;
 wire _1172_;
 wire _1173_;
 wire _1174_;
 wire _1175_;
 wire _1176_;
 wire _1177_;
 wire _1178_;
 wire _1179_;
 wire _1180_;
 wire _1181_;
 wire _1182_;
 wire _1183_;
 wire _1184_;
 wire _1185_;
 wire _1186_;
 wire _1187_;
 wire _1188_;
 wire _1189_;
 wire _1190_;
 wire _1191_;
 wire _1192_;
 wire _1193_;
 wire _1194_;
 wire _1195_;
 wire _1196_;
 wire _1197_;
 wire _1198_;
 wire _1199_;
 wire _1200_;
 wire _1201_;
 wire _1202_;
 wire _1203_;
 wire _1204_;
 wire _1205_;
 wire _1206_;
 wire _1207_;
 wire _1208_;
 wire _1209_;
 wire _1210_;
 wire _1211_;
 wire _1212_;
 wire _1213_;
 wire _1214_;
 wire _1215_;
 wire _1216_;
 wire _1217_;
 wire _1218_;
 wire _1219_;
 wire _1220_;
 wire _1221_;
 wire _1222_;
 wire _1223_;
 wire _1224_;
 wire _1225_;
 wire _1226_;
 wire _1227_;
 wire _1228_;
 wire _1229_;
 wire _1230_;
 wire _1231_;
 wire _1232_;
 wire _1233_;
 wire _1234_;
 wire _1235_;
 wire _1236_;
 wire _1237_;
 wire _1238_;
 wire _1239_;
 wire _1240_;
 wire _1241_;
 wire _1242_;
 wire _1243_;
 wire _1244_;
 wire _1245_;
 wire _1246_;
 wire _1247_;
 wire _1248_;
 wire _1249_;
 wire _1250_;
 wire _1251_;
 wire _1252_;
 wire _1253_;
 wire _1254_;
 wire _1255_;
 wire _1256_;
 wire _1257_;
 wire _1258_;
 wire _1259_;
 wire _1260_;
 wire _1261_;
 wire _1262_;
 wire _1263_;
 wire _1264_;
 wire _1265_;
 wire _1266_;
 wire _1267_;
 wire _1268_;
 wire _1269_;
 wire _1270_;
 wire _1271_;
 wire _1272_;
 wire _1273_;
 wire _1274_;
 wire _1275_;
 wire _1276_;
 wire _1277_;
 wire _1278_;
 wire _1279_;
 wire _1280_;
 wire _1281_;
 wire _1282_;
 wire _1283_;
 wire _1284_;
 wire _1285_;
 wire _1286_;
 wire _1287_;
 wire _1288_;
 wire _1289_;
 wire _1290_;
 wire _1291_;
 wire _1292_;
 wire _1293_;
 wire _1294_;
 wire _1295_;
 wire _1296_;
 wire _1297_;
 wire _1298_;
 wire _1299_;
 wire _1300_;
 wire _1301_;
 wire _1302_;
 wire _1303_;
 wire _1304_;
 wire _1305_;
 wire _1306_;
 wire _1307_;
 wire _1308_;
 wire _1309_;
 wire _1310_;
 wire _1311_;
 wire _1312_;
 wire _1313_;
 wire _1314_;
 wire _1315_;
 wire _1316_;
 wire _1317_;
 wire _1318_;
 wire _1319_;
 wire _1320_;
 wire _1321_;
 wire _1322_;
 wire _1323_;
 wire _1324_;
 wire _1325_;
 wire _1326_;
 wire _1327_;
 wire _1328_;
 wire _1329_;
 wire _1330_;
 wire _1331_;
 wire _1332_;
 wire _1333_;
 wire _1334_;
 wire _1335_;
 wire _1336_;
 wire _1337_;
 wire _1338_;
 wire _1339_;
 wire _1340_;
 wire _1341_;
 wire _1342_;
 wire _1343_;
 wire _1344_;
 wire _1345_;
 wire _1346_;
 wire _1347_;
 wire _1348_;
 wire _1349_;
 wire _1350_;
 wire _1351_;
 wire _1352_;
 wire _1353_;
 wire _1354_;
 wire _1355_;
 wire _1356_;
 wire _1357_;
 wire _1358_;
 wire _1359_;
 wire _1360_;
 wire _1361_;
 wire _1362_;
 wire _1363_;
 wire _1364_;
 wire _1365_;
 wire _1366_;
 wire _1367_;
 wire _1368_;
 wire _1369_;
 wire _1370_;
 wire _1371_;
 wire _1372_;
 wire _1373_;
 wire _1374_;
 wire _1375_;
 wire _1376_;
 wire _1377_;
 wire _1378_;
 wire _1379_;
 wire _1380_;
 wire _1381_;
 wire _1382_;
 wire _1383_;
 wire _1384_;
 wire _1385_;
 wire _1386_;
 wire _1387_;
 wire _1388_;
 wire _1389_;
 wire _1390_;
 wire _1391_;
 wire _1392_;
 wire _1393_;
 wire _1394_;
 wire _1395_;
 wire _1396_;
 wire _1397_;
 wire _1398_;
 wire _1399_;
 wire _1400_;
 wire _1401_;
 wire _1402_;
 wire _1403_;
 wire _1404_;
 wire _1405_;
 wire _1406_;
 wire _1407_;
 wire _1408_;
 wire _1409_;
 wire _1410_;
 wire _1411_;
 wire _1412_;
 wire _1413_;
 wire _1414_;
 wire _1415_;
 wire _1416_;
 wire _1417_;
 wire _1418_;
 wire _1419_;
 wire _1420_;
 wire _1421_;
 wire _1422_;
 wire _1423_;
 wire _1424_;
 wire _1425_;
 wire _1426_;
 wire _1427_;
 wire _1428_;
 wire _1429_;
 wire _1430_;
 wire _1431_;
 wire _1432_;
 wire _1433_;
 wire _1434_;
 wire _1435_;
 wire _1436_;
 wire _1437_;
 wire _1438_;
 wire _1439_;
 wire _1440_;
 wire _1441_;
 wire _1442_;
 wire _1443_;
 wire _1444_;
 wire _1445_;
 wire _1446_;
 wire _1447_;
 wire _1448_;
 wire _1449_;
 wire _1450_;
 wire _1451_;
 wire _1452_;
 wire _1453_;
 wire _1454_;
 wire _1455_;
 wire _1456_;
 wire _1457_;
 wire _1458_;
 wire _1459_;
 wire _1460_;
 wire _1461_;
 wire _1462_;
 wire _1463_;
 wire _1464_;
 wire _1465_;
 wire _1466_;
 wire _1467_;
 wire _1468_;
 wire _1469_;
 wire _1470_;
 wire _1471_;
 wire _1472_;
 wire _1473_;
 wire _1474_;
 wire _1475_;
 wire _1476_;
 wire _1477_;
 wire _1478_;
 wire _1479_;
 wire _1480_;
 wire _1481_;
 wire _1482_;
 wire _1483_;
 wire _1484_;
 wire _1485_;
 wire _1486_;
 wire _1487_;
 wire _1488_;
 wire _1489_;
 wire _1490_;
 wire _1491_;
 wire _1492_;
 wire _1493_;
 wire _1494_;
 wire _1495_;
 wire _1496_;
 wire _1497_;
 wire _1498_;
 wire _1499_;
 wire _1500_;
 wire _1501_;
 wire _1502_;
 wire _1503_;
 wire _1504_;
 wire _1505_;
 wire _1506_;
 wire _1507_;
 wire _1508_;
 wire _1509_;
 wire _1510_;
 wire _1511_;
 wire _1512_;
 wire _1513_;
 wire _1514_;
 wire _1515_;
 wire _1516_;
 wire _1517_;
 wire _1518_;
 wire _1519_;
 wire _1520_;
 wire _1521_;
 wire _1522_;
 wire _1523_;
 wire _1524_;
 wire _1525_;
 wire _1526_;
 wire _1527_;
 wire _1528_;
 wire _1529_;
 wire _1530_;
 wire _1531_;
 wire _1532_;
 wire _1533_;
 wire _1534_;
 wire _1535_;
 wire _1536_;
 wire _1537_;
 wire _1538_;
 wire _1539_;
 wire _1540_;
 wire _1541_;
 wire _1542_;
 wire _1543_;
 wire _1544_;
 wire _1545_;
 wire _1546_;
 wire _1547_;
 wire _1548_;
 wire _1549_;
 wire _1550_;
 wire _1551_;
 wire _1552_;
 wire _1553_;
 wire _1554_;
 wire _1555_;
 wire _1556_;
 wire _1557_;
 wire _1558_;
 wire _1559_;
 wire _1560_;
 wire _1561_;
 wire _1562_;
 wire _1563_;
 wire _1564_;
 wire _1565_;
 wire _1566_;
 wire _1567_;
 wire _1568_;
 wire _1569_;
 wire _1570_;
 wire _1571_;
 wire _1572_;
 wire _1573_;
 wire _1574_;
 wire _1575_;
 wire _1576_;
 wire _1577_;
 wire _1578_;
 wire _1579_;
 wire _1580_;
 wire _1581_;
 wire _1582_;
 wire _1583_;
 wire _1584_;
 wire _1585_;
 wire _1586_;
 wire _1587_;
 wire _1588_;
 wire _1589_;
 wire _1590_;
 wire _1591_;
 wire _1592_;
 wire _1593_;
 wire _1594_;
 wire _1595_;
 wire _1596_;
 wire _1597_;
 wire _1598_;
 wire _1599_;
 wire _1600_;
 wire _1601_;
 wire _1602_;
 wire _1603_;
 wire _1604_;
 wire _1605_;
 wire _1606_;
 wire _1607_;
 wire _1608_;
 wire _1609_;
 wire _1610_;
 wire _1611_;
 wire _1612_;
 wire _1613_;
 wire _1614_;
 wire _1615_;
 wire _1616_;
 wire _1617_;
 wire _1618_;
 wire _1619_;
 wire _1620_;
 wire _1621_;
 wire _1622_;
 wire _1623_;
 wire _1624_;
 wire _1625_;
 wire _1626_;
 wire _1627_;
 wire _1628_;
 wire _1629_;
 wire _1630_;
 wire _1631_;
 wire _1632_;
 wire _1633_;
 wire _1634_;
 wire _1635_;
 wire _1636_;
 wire _1637_;
 wire _1638_;
 wire _1639_;
 wire _1640_;
 wire _1641_;
 wire _1642_;
 wire _1643_;
 wire _1644_;
 wire _1645_;
 wire _1646_;
 wire _1647_;
 wire _1648_;
 wire _1649_;
 wire _1650_;
 wire _1651_;
 wire _1652_;
 wire _1653_;
 wire _1654_;
 wire _1655_;
 wire _1656_;
 wire _1657_;
 wire _1658_;
 wire _1659_;
 wire _1660_;
 wire _1661_;
 wire _1662_;
 wire _1663_;
 wire _1664_;
 wire _1665_;
 wire _1666_;
 wire _1667_;
 wire _1668_;
 wire _1669_;
 wire _1670_;
 wire _1671_;
 wire _1672_;
 wire _1673_;
 wire _1674_;
 wire _1675_;
 wire _1676_;
 wire _1677_;
 wire _1678_;
 wire _1679_;
 wire _1680_;
 wire _1681_;
 wire _1682_;
 wire _1683_;
 wire _1684_;
 wire _1685_;
 wire _1686_;
 wire _1687_;
 wire _1688_;
 wire _1689_;
 wire _1690_;
 wire _1691_;
 wire _1692_;
 wire _1693_;
 wire _1694_;
 wire _1695_;
 wire _1696_;
 wire _1697_;
 wire _1698_;
 wire _1699_;
 wire _1700_;
 wire _1701_;
 wire _1702_;
 wire _1703_;
 wire _1704_;
 wire _1705_;
 wire _1706_;
 wire _1707_;
 wire _1708_;
 wire _1709_;
 wire _1710_;
 wire _1711_;
 wire _1712_;
 wire _1713_;
 wire _1714_;
 wire _1715_;
 wire _1716_;
 wire _1717_;
 wire _1718_;
 wire _1719_;
 wire _1720_;
 wire _1721_;
 wire _1722_;
 wire _1723_;
 wire _1724_;
 wire _1725_;
 wire _1726_;
 wire _1727_;
 wire _1728_;
 wire _1729_;
 wire _1730_;
 wire _1731_;
 wire _1732_;
 wire _1733_;
 wire _1734_;
 wire _1735_;
 wire _1736_;
 wire _1737_;
 wire _1738_;
 wire _1739_;
 wire _1740_;
 wire _1741_;
 wire _1742_;
 wire _1743_;
 wire _1744_;
 wire _1745_;
 wire _1746_;
 wire _1747_;
 wire _1748_;
 wire _1749_;
 wire _1750_;
 wire _1751_;
 wire _1752_;
 wire _1753_;
 wire _1754_;
 wire _1755_;
 wire _1756_;
 wire _1757_;
 wire _1758_;
 wire _1759_;
 wire _1760_;
 wire _1761_;
 wire _1762_;
 wire _1763_;
 wire _1764_;
 wire _1765_;
 wire _1766_;
 wire _1767_;
 wire _1768_;
 wire _1769_;
 wire _1770_;
 wire _1771_;
 wire _1772_;
 wire _1773_;
 wire _1774_;
 wire _1775_;
 wire _1776_;
 wire _1777_;
 wire _1778_;
 wire _1779_;
 wire _1780_;
 wire _1781_;
 wire _1782_;
 wire _1783_;
 wire _1784_;
 wire _1785_;
 wire _1786_;
 wire _1787_;
 wire _1788_;
 wire _1789_;
 wire _1790_;
 wire _1791_;
 wire _1792_;
 wire _1793_;
 wire _1794_;
 wire _1795_;
 wire _1796_;
 wire _1797_;
 wire _1798_;
 wire _1799_;
 wire _1800_;
 wire _1801_;
 wire _1802_;
 wire _1803_;
 wire _1804_;
 wire _1805_;
 wire _1806_;
 wire _1807_;
 wire _1808_;
 wire _1809_;
 wire _1810_;
 wire _1811_;
 wire _1812_;
 wire _1813_;
 wire _1814_;
 wire _1815_;
 wire _1816_;
 wire _1817_;
 wire _1818_;
 wire _1819_;
 wire _1820_;
 wire _1821_;
 wire _1822_;
 wire _1823_;
 wire _1824_;
 wire _1825_;
 wire _1826_;
 wire _1827_;
 wire _1828_;
 wire _1829_;
 wire _1830_;
 wire _1831_;
 wire _1832_;
 wire _1833_;
 wire _1834_;
 wire _1835_;
 wire _1836_;
 wire _1837_;
 wire _1838_;
 wire _1839_;
 wire _1840_;
 wire _1841_;
 wire _1842_;
 wire _1843_;
 wire _1844_;
 wire _1845_;
 wire _1846_;
 wire _1847_;
 wire _1848_;
 wire _1849_;
 wire _1850_;
 wire _1851_;
 wire _1852_;
 wire _1853_;
 wire _1854_;
 wire _1855_;
 wire _1856_;
 wire _1857_;
 wire _1858_;
 wire _1859_;
 wire _1860_;
 wire _1861_;
 wire _1862_;
 wire _1863_;
 wire _1864_;
 wire _1865_;
 wire _1866_;
 wire _1867_;
 wire _1868_;
 wire _1869_;
 wire _1870_;
 wire _1871_;
 wire _1872_;
 wire _1873_;
 wire _1874_;
 wire _1875_;
 wire _1876_;
 wire _1877_;
 wire _1878_;
 wire _1879_;
 wire _1880_;
 wire _1881_;
 wire _1882_;
 wire _1883_;
 wire _1884_;
 wire _1885_;
 wire _1886_;
 wire _1887_;
 wire _1888_;
 wire _1889_;
 wire _1890_;
 wire _1891_;
 wire _1892_;
 wire _1893_;
 wire _1894_;
 wire _1895_;
 wire _1896_;
 wire _1897_;
 wire _1898_;
 wire _1899_;
 wire _1900_;
 wire _1901_;
 wire _1902_;
 wire _1903_;
 wire _1904_;
 wire _1905_;
 wire _1906_;
 wire _1907_;
 wire _1908_;
 wire _1909_;
 wire _1910_;
 wire _1911_;
 wire _1912_;
 wire _1913_;
 wire _1914_;
 wire _1915_;
 wire _1916_;
 wire _1917_;
 wire _1918_;
 wire _1919_;
 wire _1920_;
 wire _1921_;
 wire _1922_;
 wire _1923_;
 wire _1924_;
 wire _1925_;
 wire _1926_;
 wire _1927_;
 wire _1928_;
 wire _1929_;
 wire _1930_;
 wire _1931_;
 wire _1932_;
 wire _1933_;
 wire _1934_;
 wire _1935_;
 wire _1936_;
 wire _1937_;
 wire _1938_;
 wire _1939_;
 wire _1940_;
 wire _1941_;
 wire _1942_;
 wire _1943_;
 wire _1944_;
 wire _1945_;
 wire _1946_;
 wire _1947_;
 wire _1948_;
 wire _1949_;
 wire _1950_;
 wire _1951_;
 wire _1952_;
 wire _1953_;
 wire _1954_;
 wire _1955_;
 wire _1956_;
 wire _1957_;
 wire _1958_;
 wire _1959_;
 wire _1960_;
 wire _1961_;
 wire _1962_;
 wire _1963_;
 wire _1964_;
 wire _1965_;
 wire _1966_;
 wire _1967_;
 wire _1968_;
 wire _1969_;
 wire _1970_;
 wire _1971_;
 wire _1972_;
 wire _1973_;
 wire _1974_;
 wire _1975_;
 wire _1976_;
 wire _1977_;
 wire _1978_;
 wire _1979_;
 wire _1980_;
 wire _1981_;
 wire _1982_;
 wire _1983_;
 wire _1984_;
 wire _1985_;
 wire _1986_;
 wire _1987_;
 wire _1988_;
 wire _1989_;
 wire _1990_;
 wire _1991_;
 wire _1992_;
 wire _1993_;
 wire _1994_;
 wire _1995_;
 wire _1996_;
 wire _1997_;
 wire _1998_;
 wire _1999_;
 wire _2000_;
 wire _2001_;
 wire _2002_;
 wire _2003_;
 wire _2004_;
 wire _2005_;
 wire _2006_;
 wire _2007_;
 wire _2008_;
 wire _2009_;
 wire _2010_;
 wire _2011_;
 wire _2012_;
 wire _2013_;
 wire _2014_;
 wire _2015_;
 wire _2016_;
 wire _2017_;
 wire _2018_;
 wire _2019_;
 wire _2020_;
 wire _2021_;
 wire _2022_;
 wire _2023_;
 wire _2024_;
 wire _2025_;
 wire _2026_;
 wire _2027_;
 wire _2028_;
 wire _2029_;
 wire _2030_;
 wire _2031_;
 wire _2032_;
 wire _2033_;
 wire _2034_;
 wire _2035_;
 wire _2036_;
 wire _2037_;
 wire _2038_;
 wire _2039_;
 wire _2040_;
 wire _2041_;
 wire _2042_;
 wire _2043_;
 wire _2044_;
 wire _2045_;
 wire _2046_;
 wire _2047_;
 wire _2048_;
 wire _2049_;
 wire _2050_;
 wire _2051_;
 wire _2052_;
 wire _2053_;
 wire _2054_;
 wire _2055_;
 wire _2056_;
 wire _2057_;
 wire _2058_;
 wire _2059_;
 wire _2060_;
 wire _2061_;
 wire _2062_;
 wire _2063_;
 wire _2064_;
 wire _2065_;
 wire _2066_;
 wire _2067_;
 wire _2068_;
 wire _2069_;
 wire _2070_;
 wire _2071_;
 wire _2072_;
 wire _2073_;
 wire _2074_;
 wire _2075_;
 wire _2076_;
 wire _2077_;
 wire _2078_;
 wire _2079_;
 wire _2080_;
 wire _2081_;
 wire _2082_;
 wire _2083_;
 wire _2084_;
 wire _2085_;
 wire _2086_;
 wire _2087_;
 wire _2088_;
 wire _2089_;
 wire _2090_;
 wire _2091_;
 wire _2092_;
 wire _2093_;
 wire _2094_;
 wire _2095_;
 wire _2096_;
 wire _2097_;
 wire _2098_;
 wire _2099_;
 wire _2100_;
 wire _2101_;
 wire _2102_;
 wire _2103_;
 wire _2104_;
 wire _2105_;
 wire _2106_;
 wire _2107_;
 wire _2108_;
 wire _2109_;
 wire _2110_;
 wire _2111_;
 wire _2112_;
 wire _2113_;
 wire _2114_;
 wire _2115_;
 wire _2116_;
 wire _2117_;
 wire _2118_;
 wire _2119_;
 wire _2120_;
 wire _2121_;
 wire _2122_;
 wire _2123_;
 wire _2124_;
 wire _2125_;
 wire _2126_;
 wire _2127_;
 wire _2128_;
 wire _2129_;
 wire _2130_;
 wire _2131_;
 wire _2132_;
 wire _2133_;
 wire _2134_;
 wire _2135_;
 wire _2136_;
 wire _2137_;
 wire _2138_;
 wire _2139_;
 wire _2140_;
 wire _2141_;
 wire _2142_;
 wire _2143_;
 wire _2144_;
 wire _2145_;
 wire _2146_;
 wire _2147_;
 wire _2148_;
 wire _2149_;
 wire _2150_;
 wire _2151_;
 wire _2152_;
 wire _2153_;
 wire _2154_;
 wire _2155_;
 wire _2156_;
 wire _2157_;
 wire _2158_;
 wire _2159_;
 wire _2160_;
 wire _2161_;
 wire _2162_;
 wire _2163_;
 wire _2164_;
 wire _2165_;
 wire _2166_;
 wire _2167_;
 wire _2168_;
 wire _2169_;
 wire _2170_;
 wire _2171_;
 wire _2172_;
 wire _2173_;
 wire _2174_;
 wire _2175_;
 wire _2176_;
 wire _2177_;
 wire _2178_;
 wire _2179_;
 wire _2180_;
 wire _2181_;
 wire _2182_;
 wire _2183_;
 wire _2184_;
 wire _2185_;
 wire _2186_;
 wire _2187_;
 wire _2188_;
 wire _2189_;
 wire _2190_;
 wire _2191_;
 wire _2192_;
 wire _2193_;
 wire _2194_;
 wire _2195_;
 wire _2196_;
 wire _2197_;
 wire _2198_;
 wire _2199_;
 wire _2200_;
 wire _2201_;
 wire _2202_;
 wire _2203_;
 wire _2204_;
 wire _2205_;
 wire _2206_;
 wire _2207_;
 wire _2208_;
 wire _2209_;
 wire _2210_;
 wire _2211_;
 wire _2212_;
 wire _2213_;
 wire _2214_;
 wire _2215_;
 wire _2216_;
 wire _2217_;
 wire _2218_;
 wire _2219_;
 wire _2220_;
 wire _2221_;
 wire _2222_;
 wire _2223_;
 wire _2224_;
 wire _2225_;
 wire _2226_;
 wire _2227_;
 wire _2228_;
 wire _2229_;
 wire _2230_;
 wire _2231_;
 wire _2232_;
 wire _2233_;
 wire _2234_;
 wire _2235_;
 wire _2236_;
 wire _2237_;
 wire _2238_;
 wire _2239_;
 wire _2240_;
 wire _2241_;
 wire _2242_;
 wire _2243_;
 wire _2244_;
 wire _2245_;
 wire _2246_;
 wire _2247_;
 wire _2248_;
 wire _2249_;
 wire _2250_;
 wire _2251_;
 wire _2252_;
 wire _2253_;
 wire _2254_;
 wire _2255_;
 wire _2256_;
 wire _2257_;
 wire _2258_;
 wire _2259_;
 wire _2260_;
 wire _2261_;
 wire _2262_;
 wire _2263_;
 wire _2264_;
 wire _2265_;
 wire _2266_;
 wire _2267_;
 wire _2268_;
 wire _2269_;
 wire _2270_;
 wire _2271_;
 wire _2272_;
 wire _2273_;
 wire _2274_;
 wire _2275_;
 wire _2276_;
 wire _2277_;
 wire _2278_;
 wire _2279_;
 wire _2280_;
 wire _2281_;
 wire _2282_;
 wire _2283_;
 wire _2284_;
 wire _2285_;
 wire _2286_;
 wire _2287_;
 wire _2288_;
 wire _2289_;
 wire _2290_;
 wire _2291_;
 wire _2292_;
 wire _2293_;
 wire _2294_;
 wire _2295_;
 wire _2296_;
 wire _2297_;
 wire _2298_;
 wire _2299_;
 wire _2300_;
 wire _2301_;
 wire _2302_;
 wire _2303_;
 wire _2304_;
 wire _2305_;
 wire _2306_;
 wire _2307_;
 wire _2308_;
 wire _2309_;
 wire _2310_;
 wire _2311_;
 wire _2312_;
 wire _2313_;
 wire _2314_;
 wire _2315_;
 wire _2316_;
 wire _2317_;
 wire _2318_;
 wire _2319_;
 wire _2320_;
 wire _2321_;
 wire _2322_;
 wire _2323_;
 wire _2324_;
 wire _2325_;
 wire _2326_;
 wire _2327_;
 wire _2328_;
 wire _2329_;
 wire _2330_;
 wire _2331_;
 wire _2332_;
 wire _2333_;
 wire _2334_;
 wire _2335_;
 wire _2336_;
 wire _2337_;
 wire _2338_;
 wire _2339_;
 wire _2340_;
 wire _2341_;
 wire _2342_;
 wire _2343_;
 wire _2344_;
 wire _2345_;
 wire _2346_;
 wire _2347_;
 wire _2348_;
 wire _2349_;
 wire _2350_;
 wire _2351_;
 wire _2352_;
 wire _2353_;
 wire _2354_;
 wire _2355_;
 wire _2356_;
 wire _2357_;
 wire _2358_;
 wire _2359_;
 wire _2360_;
 wire _2361_;
 wire _2362_;
 wire _2363_;
 wire _2364_;
 wire _2365_;
 wire _2366_;
 wire _2367_;
 wire _2368_;
 wire _2369_;
 wire _2370_;
 wire _2371_;
 wire _2372_;
 wire _2373_;
 wire _2374_;
 wire _2375_;
 wire _2376_;
 wire _2377_;
 wire _2378_;
 wire _2379_;
 wire _2380_;
 wire _2381_;
 wire _2382_;
 wire _2383_;
 wire _2384_;
 wire _2385_;
 wire _2386_;
 wire _2387_;
 wire _2388_;
 wire _2389_;
 wire _2390_;
 wire _2391_;
 wire _2392_;
 wire _2393_;
 wire _2394_;
 wire _2395_;
 wire _2396_;
 wire _2397_;
 wire _2398_;
 wire _2399_;
 wire _2400_;
 wire _2401_;
 wire _2402_;
 wire _2403_;
 wire _2404_;
 wire _2405_;
 wire _2406_;
 wire _2407_;
 wire _2408_;
 wire _2409_;
 wire _2410_;
 wire _2411_;
 wire _2412_;
 wire _2413_;
 wire _2414_;
 wire _2415_;
 wire _2416_;
 wire _2417_;
 wire _2418_;
 wire _2419_;
 wire _2420_;
 wire _2421_;
 wire _2422_;
 wire _2423_;
 wire _2424_;
 wire _2425_;
 wire _2426_;
 wire _2427_;
 wire _2428_;
 wire _2429_;
 wire _2430_;
 wire _2431_;
 wire _2432_;
 wire _2433_;
 wire _2434_;
 wire _2435_;
 wire _2436_;
 wire _2437_;
 wire _2438_;
 wire _2439_;
 wire _2440_;
 wire _2441_;
 wire _2442_;
 wire _2443_;
 wire _2444_;
 wire _2445_;
 wire _2446_;
 wire _2447_;
 wire _2448_;
 wire _2449_;
 wire _2450_;
 wire _2451_;
 wire _2452_;
 wire _2453_;
 wire _2454_;
 wire _2455_;
 wire _2456_;
 wire _2457_;
 wire _2458_;
 wire _2459_;
 wire _2460_;
 wire _2461_;
 wire _2462_;
 wire _2463_;
 wire _2464_;
 wire _2465_;
 wire _2466_;
 wire _2467_;
 wire _2468_;
 wire _2469_;
 wire _2470_;
 wire _2471_;
 wire _2472_;
 wire _2473_;
 wire _2474_;
 wire _2475_;
 wire _2476_;
 wire _2477_;
 wire _2478_;
 wire _2479_;
 wire _2480_;
 wire _2481_;
 wire _2482_;
 wire _2483_;
 wire _2484_;
 wire _2485_;
 wire _2486_;
 wire _2487_;
 wire _2488_;
 wire _2489_;
 wire _2490_;
 wire _2491_;
 wire _2492_;
 wire _2493_;
 wire _2494_;
 wire _2495_;
 wire _2496_;
 wire _2497_;
 wire _2498_;
 wire _2499_;
 wire _2500_;
 wire _2501_;
 wire _2502_;
 wire _2503_;
 wire _2504_;
 wire _2505_;
 wire _2506_;
 wire _2507_;
 wire _2508_;
 wire _2509_;
 wire _2510_;
 wire _2511_;
 wire _2512_;
 wire _2513_;
 wire _2514_;
 wire _2515_;
 wire _2516_;
 wire _2517_;
 wire _2518_;
 wire _2519_;
 wire _2520_;
 wire _2521_;
 wire _2522_;
 wire _2523_;
 wire _2524_;
 wire _2525_;
 wire _2526_;
 wire _2527_;
 wire _2528_;
 wire _2529_;
 wire _2530_;
 wire _2531_;
 wire _2532_;
 wire _2533_;
 wire _2534_;
 wire _2535_;
 wire _2536_;
 wire _2537_;
 wire _2538_;
 wire _2539_;
 wire _2540_;
 wire _2541_;
 wire _2542_;
 wire _2543_;
 wire _2544_;
 wire _2545_;
 wire _2546_;
 wire _2547_;
 wire _2548_;
 wire _2549_;
 wire _2550_;
 wire _2551_;
 wire _2552_;
 wire _2553_;
 wire _2554_;
 wire _2555_;
 wire _2556_;
 wire _2557_;
 wire _2558_;
 wire _2559_;
 wire _2560_;
 wire _2561_;
 wire _2562_;
 wire _2563_;
 wire _2564_;
 wire _2565_;
 wire _2566_;
 wire _2567_;
 wire _2568_;
 wire _2569_;
 wire _2570_;
 wire _2571_;
 wire _2572_;
 wire _2573_;
 wire _2574_;
 wire _2575_;
 wire _2576_;
 wire _2577_;
 wire _2578_;
 wire _2579_;
 wire _2580_;
 wire _2581_;
 wire _2582_;
 wire _2583_;
 wire _2584_;
 wire _2585_;
 wire _2586_;
 wire _2587_;
 wire _2588_;
 wire _2589_;
 wire _2590_;
 wire _2591_;
 wire _2592_;
 wire _2593_;
 wire _2594_;
 wire _2595_;
 wire _2596_;
 wire _2597_;
 wire _2598_;
 wire _2599_;
 wire _2600_;
 wire _2601_;
 wire _2602_;
 wire _2603_;
 wire _2604_;
 wire _2605_;
 wire _2606_;
 wire _2607_;
 wire _2608_;
 wire _2609_;
 wire _2610_;
 wire _2611_;
 wire _2612_;
 wire _2613_;
 wire _2614_;
 wire _2615_;
 wire _2616_;
 wire _2617_;
 wire _2618_;
 wire _2619_;
 wire _2620_;
 wire _2621_;
 wire _2622_;
 wire _2623_;
 wire _2624_;
 wire _2625_;
 wire _2626_;
 wire _2627_;
 wire _2628_;
 wire _2629_;
 wire _2630_;
 wire _2631_;
 wire _2632_;
 wire _2633_;
 wire _2634_;
 wire _2635_;
 wire _2636_;
 wire _2637_;
 wire _2638_;
 wire _2639_;
 wire _2640_;
 wire _2641_;
 wire _2642_;
 wire _2643_;
 wire _2644_;
 wire _2645_;
 wire _2646_;
 wire _2647_;
 wire _2648_;
 wire _2649_;
 wire _2650_;
 wire _2651_;
 wire _2652_;
 wire _2653_;
 wire _2654_;
 wire _2655_;
 wire _2656_;
 wire _2657_;
 wire _2658_;
 wire _2659_;
 wire _2660_;
 wire _2661_;
 wire _2662_;
 wire _2663_;
 wire _2664_;
 wire _2665_;
 wire _2666_;
 wire _2667_;
 wire _2668_;
 wire _2669_;
 wire _2670_;
 wire _2671_;
 wire _2672_;
 wire _2673_;
 wire _2674_;
 wire _2675_;
 wire _2676_;
 wire _2677_;
 wire _2678_;
 wire _2679_;
 wire _2680_;
 wire _2681_;
 wire _2682_;
 wire _2683_;
 wire _2684_;
 wire _2685_;
 wire _2686_;
 wire _2687_;
 wire _2688_;
 wire _2689_;
 wire _2690_;
 wire _2691_;
 wire _2692_;
 wire _2693_;
 wire _2694_;
 wire _2695_;
 wire _2696_;
 wire _2697_;
 wire _2698_;
 wire _2699_;
 wire _2700_;
 wire _2701_;
 wire _2702_;
 wire _2703_;
 wire _2704_;
 wire _2705_;
 wire _2706_;
 wire _2707_;
 wire _2708_;
 wire _2709_;
 wire _2710_;
 wire _2711_;
 wire _2712_;
 wire _2713_;
 wire _2714_;
 wire _2715_;
 wire _2716_;
 wire _2717_;
 wire _2718_;
 wire _2719_;
 wire _2720_;
 wire _2721_;
 wire _2722_;
 wire _2723_;
 wire _2724_;
 wire _2725_;
 wire _2726_;
 wire _2727_;
 wire _2728_;
 wire _2729_;
 wire _2730_;
 wire _2731_;
 wire _2732_;
 wire _2733_;
 wire _2734_;
 wire _2735_;
 wire _2736_;
 wire _2737_;
 wire _2738_;
 wire _2739_;
 wire _2740_;
 wire _2741_;
 wire _2742_;
 wire _2743_;
 wire _2744_;
 wire _2745_;
 wire _2746_;
 wire _2747_;
 wire _2748_;
 wire _2749_;
 wire _2750_;
 wire _2751_;
 wire _2752_;
 wire _2753_;
 wire _2754_;
 wire _2755_;
 wire _2756_;
 wire _2757_;
 wire _2758_;
 wire _2759_;
 wire _2760_;
 wire _2761_;
 wire _2762_;
 wire _2763_;
 wire _2764_;
 wire _2765_;
 wire _2766_;
 wire _2767_;
 wire _2768_;
 wire _2769_;
 wire _2770_;
 wire _2771_;
 wire _2772_;
 wire _2773_;
 wire _2774_;
 wire _2775_;
 wire _2776_;
 wire _2777_;
 wire _2778_;
 wire _2779_;
 wire _2780_;
 wire _2781_;
 wire _2782_;
 wire _2783_;
 wire _2784_;
 wire _2785_;
 wire _2786_;
 wire _2787_;
 wire _2788_;
 wire _2789_;
 wire _2790_;
 wire _2791_;
 wire _2792_;
 wire _2793_;
 wire _2794_;
 wire _2795_;
 wire _2796_;
 wire _2797_;
 wire _2798_;
 wire _2799_;
 wire _2800_;
 wire _2801_;
 wire _2802_;
 wire _2803_;
 wire _2804_;
 wire _2805_;
 wire _2806_;
 wire _2807_;
 wire _2808_;
 wire _2809_;
 wire _2810_;
 wire _2811_;
 wire _2812_;
 wire _2813_;
 wire _2814_;
 wire _2815_;
 wire _2816_;
 wire _2817_;
 wire _2818_;
 wire _2819_;
 wire _2820_;
 wire _2821_;
 wire _2822_;
 wire _2823_;
 wire _2824_;
 wire _2825_;
 wire _2826_;
 wire _2827_;
 wire _2828_;
 wire _2829_;
 wire _2830_;
 wire _2831_;
 wire _2832_;
 wire _2833_;
 wire _2834_;
 wire _2835_;
 wire _2836_;
 wire _2837_;
 wire _2838_;
 wire _2839_;
 wire _2840_;
 wire _2841_;
 wire _2842_;
 wire _2843_;
 wire _2844_;
 wire _2845_;
 wire _2846_;
 wire _2847_;
 wire _2848_;
 wire _2849_;
 wire _2850_;
 wire _2851_;
 wire _2852_;
 wire _2853_;
 wire _2854_;
 wire _2855_;
 wire _2856_;
 wire _2857_;
 wire _2858_;
 wire _2859_;
 wire _2860_;
 wire _2861_;
 wire _2862_;
 wire _2863_;
 wire _2864_;
 wire _2865_;
 wire _2866_;
 wire _2867_;
 wire _2868_;
 wire _2869_;
 wire _2870_;
 wire _2871_;
 wire _2872_;
 wire _2873_;
 wire _2874_;
 wire _2875_;
 wire _2876_;
 wire _2877_;
 wire _2878_;
 wire _2879_;
 wire _2880_;
 wire _2881_;
 wire _2882_;
 wire _2883_;
 wire _2884_;
 wire _2885_;
 wire _2886_;
 wire _2887_;
 wire _2888_;
 wire _2889_;
 wire _2890_;
 wire _2891_;
 wire _2892_;
 wire _2893_;
 wire _2894_;
 wire _2895_;
 wire _2896_;
 wire _2897_;
 wire _2898_;
 wire _2899_;
 wire _2900_;
 wire _2901_;
 wire _2902_;
 wire _2903_;
 wire _2904_;
 wire _2905_;
 wire _2906_;
 wire _2907_;
 wire _2908_;
 wire _2909_;
 wire _2910_;
 wire _2911_;
 wire _2912_;
 wire _2913_;
 wire _2914_;
 wire _2915_;
 wire _2916_;
 wire _2917_;
 wire _2918_;
 wire _2919_;
 wire _2920_;
 wire _2921_;
 wire _2922_;
 wire _2923_;
 wire _2924_;
 wire _2925_;
 wire _2926_;
 wire _2927_;
 wire _2928_;
 wire _2929_;
 wire _2930_;
 wire _2931_;
 wire _2932_;
 wire _2933_;
 wire _2934_;
 wire _2935_;
 wire _2936_;
 wire _2937_;
 wire _2938_;
 wire _2939_;
 wire _2940_;
 wire _2941_;
 wire _2942_;
 wire _2943_;
 wire _2944_;
 wire _2945_;
 wire _2946_;
 wire _2947_;
 wire _2948_;
 wire _2949_;
 wire _2950_;
 wire _2951_;
 wire _2952_;
 wire _2953_;
 wire _2954_;
 wire _2955_;
 wire _2956_;
 wire _2957_;
 wire _2958_;
 wire _2959_;
 wire _2960_;
 wire _2961_;
 wire _2962_;
 wire _2963_;
 wire _2964_;
 wire _2965_;
 wire _2966_;
 wire _2967_;
 wire _2968_;
 wire _2969_;
 wire _2970_;
 wire _2971_;
 wire _2972_;
 wire _2973_;
 wire _2974_;
 wire _2975_;
 wire _2976_;
 wire _2977_;
 wire _2978_;
 wire _2979_;
 wire _2980_;
 wire _2981_;
 wire _2982_;
 wire _2983_;
 wire _2984_;
 wire _2985_;
 wire _2986_;
 wire _2987_;
 wire _2988_;
 wire _2989_;
 wire _2990_;
 wire _2991_;
 wire _2992_;
 wire _2993_;
 wire _2994_;
 wire _2995_;
 wire _2996_;
 wire _2997_;
 wire _2998_;
 wire _2999_;
 wire _3000_;
 wire _3001_;
 wire _3002_;
 wire _3003_;
 wire _3004_;
 wire _3005_;
 wire _3006_;
 wire _3007_;
 wire _3008_;
 wire _3009_;
 wire _3010_;
 wire _3011_;
 wire _3012_;
 wire _3013_;
 wire _3014_;
 wire _3015_;
 wire _3016_;
 wire _3017_;
 wire _3018_;
 wire _3019_;
 wire _3020_;
 wire _3021_;
 wire _3022_;
 wire _3023_;
 wire _3024_;
 wire _3025_;
 wire _3026_;
 wire _3027_;
 wire _3028_;
 wire _3029_;
 wire _3030_;
 wire _3031_;
 wire _3032_;
 wire _3033_;
 wire _3034_;
 wire _3035_;
 wire _3036_;
 wire _3037_;
 wire _3038_;
 wire _3039_;
 wire _3040_;
 wire _3041_;
 wire _3042_;
 wire _3043_;
 wire _3044_;
 wire _3045_;
 wire _3046_;
 wire _3047_;
 wire _3048_;
 wire _3049_;
 wire _3050_;
 wire _3051_;
 wire _3052_;
 wire _3053_;
 wire _3054_;
 wire _3055_;
 wire _3056_;
 wire _3057_;
 wire _3058_;
 wire _3059_;
 wire _3060_;
 wire _3061_;
 wire _3062_;
 wire _3063_;
 wire _3064_;
 wire _3065_;
 wire _3066_;
 wire _3067_;
 wire _3068_;
 wire _3069_;
 wire _3070_;
 wire _3071_;
 wire _3072_;
 wire _3073_;
 wire _3074_;
 wire _3075_;
 wire _3076_;
 wire _3077_;
 wire _3078_;
 wire _3079_;
 wire _3080_;
 wire _3081_;
 wire _3082_;
 wire _3083_;
 wire _3084_;
 wire _3085_;
 wire _3086_;
 wire _3087_;
 wire _3088_;
 wire _3089_;
 wire _3090_;
 wire _3091_;
 wire _3092_;
 wire _3093_;
 wire _3094_;
 wire _3095_;
 wire _3096_;
 wire _3097_;
 wire _3098_;
 wire _3099_;
 wire _3100_;
 wire _3101_;
 wire _3102_;
 wire _3103_;
 wire _3104_;
 wire _3105_;
 wire _3106_;
 wire _3107_;
 wire _3108_;
 wire _3109_;
 wire _3110_;
 wire _3111_;
 wire _3112_;
 wire _3113_;
 wire _3114_;
 wire _3115_;
 wire _3116_;
 wire _3117_;
 wire _3118_;
 wire _3119_;
 wire _3120_;
 wire _3121_;
 wire _3122_;
 wire _3123_;
 wire _3124_;
 wire _3125_;
 wire _3126_;
 wire _3127_;
 wire _3128_;
 wire _3129_;
 wire _3130_;
 wire _3131_;
 wire _3132_;
 wire _3133_;
 wire _3134_;
 wire _3135_;
 wire _3136_;
 wire _3137_;
 wire _3138_;
 wire _3139_;
 wire _3140_;
 wire _3141_;
 wire _3142_;
 wire _3143_;
 wire _3144_;
 wire _3145_;
 wire _3146_;
 wire _3147_;
 wire _3148_;
 wire _3149_;
 wire _3150_;
 wire _3151_;
 wire _3152_;
 wire _3153_;
 wire _3154_;
 wire _3155_;
 wire _3156_;
 wire _3157_;
 wire _3158_;
 wire _3159_;
 wire _3160_;
 wire _3161_;
 wire _3162_;
 wire _3163_;
 wire _3164_;
 wire _3165_;
 wire _3166_;
 wire _3167_;
 wire _3168_;
 wire _3169_;
 wire _3170_;
 wire _3171_;
 wire _3172_;
 wire _3173_;
 wire _3174_;
 wire _3175_;
 wire _3176_;
 wire _3177_;
 wire _3178_;
 wire _3179_;
 wire _3180_;
 wire _3181_;
 wire _3182_;
 wire _3183_;
 wire _3184_;
 wire _3185_;
 wire _3186_;
 wire _3187_;
 wire _3188_;
 wire _3189_;
 wire _3190_;
 wire _3191_;
 wire _3192_;
 wire _3193_;
 wire _3194_;
 wire _3195_;
 wire _3196_;
 wire _3197_;
 wire _3198_;
 wire _3199_;
 wire _3200_;
 wire _3201_;
 wire _3202_;
 wire _3203_;
 wire _3204_;
 wire _3205_;
 wire _3206_;
 wire _3207_;
 wire _3208_;
 wire _3209_;
 wire _3210_;
 wire _3211_;
 wire _3212_;
 wire _3213_;
 wire _3214_;
 wire _3215_;
 wire _3216_;
 wire _3217_;
 wire _3218_;
 wire _3219_;
 wire _3220_;
 wire _3221_;
 wire _3222_;
 wire _3223_;
 wire _3224_;
 wire _3225_;
 wire _3226_;
 wire _3227_;
 wire _3228_;
 wire _3229_;
 wire _3230_;
 wire _3231_;
 wire _3232_;
 wire _3233_;
 wire _3234_;
 wire _3235_;
 wire _3236_;
 wire _3237_;
 wire _3238_;
 wire _3239_;
 wire _3240_;
 wire _3241_;
 wire _3242_;
 wire _3243_;
 wire _3244_;
 wire _3245_;
 wire _3246_;
 wire _3247_;
 wire _3248_;
 wire _3249_;
 wire _3250_;
 wire _3251_;
 wire _3252_;
 wire _3253_;
 wire _3254_;
 wire _3255_;
 wire _3256_;
 wire _3257_;
 wire _3258_;
 wire _3259_;
 wire _3260_;
 wire _3261_;
 wire _3262_;
 wire _3263_;
 wire _3264_;
 wire _3265_;
 wire _3266_;
 wire _3267_;
 wire _3268_;
 wire _3269_;
 wire _3270_;
 wire _3271_;
 wire _3272_;
 wire _3273_;
 wire _3274_;
 wire _3275_;
 wire _3276_;
 wire _3277_;
 wire _3278_;
 wire _3279_;
 wire _3280_;
 wire _3281_;
 wire _3282_;
 wire _3283_;
 wire _3284_;
 wire _3285_;
 wire _3286_;
 wire _3287_;
 wire _3288_;
 wire _3289_;
 wire _3290_;
 wire _3291_;
 wire _3292_;
 wire _3293_;
 wire _3294_;
 wire _3295_;
 wire _3296_;
 wire _3297_;
 wire _3298_;
 wire _3299_;
 wire _3300_;
 wire _3301_;
 wire _3302_;
 wire _3303_;
 wire _3304_;
 wire _3305_;
 wire _3306_;
 wire _3307_;
 wire _3308_;
 wire _3309_;
 wire _3310_;
 wire _3311_;
 wire _3312_;
 wire _3313_;
 wire _3314_;
 wire _3315_;
 wire _3316_;
 wire _3317_;
 wire _3318_;
 wire _3319_;
 wire _3320_;
 wire _3321_;
 wire _3322_;
 wire _3323_;
 wire _3324_;
 wire _3325_;
 wire _3326_;
 wire _3327_;
 wire _3328_;
 wire _3329_;
 wire _3330_;
 wire _3331_;
 wire _3332_;
 wire _3333_;
 wire _3334_;
 wire _3335_;
 wire _3336_;
 wire _3337_;
 wire _3338_;
 wire _3339_;
 wire _3340_;
 wire _3341_;
 wire _3342_;
 wire _3343_;
 wire _3344_;
 wire _3345_;
 wire _3346_;
 wire _3347_;
 wire _3348_;
 wire _3349_;
 wire _3350_;
 wire _3351_;
 wire _3352_;
 wire _3353_;
 wire _3354_;
 wire _3355_;
 wire _3356_;
 wire _3357_;
 wire _3358_;
 wire _3359_;
 wire _3360_;
 wire _3361_;
 wire _3362_;
 wire _3363_;
 wire _3364_;
 wire _3365_;
 wire _3366_;
 wire _3367_;
 wire _3368_;
 wire _3369_;
 wire _3370_;
 wire _3371_;
 wire _3372_;
 wire _3373_;
 wire _3374_;
 wire _3375_;
 wire _3376_;
 wire _3377_;
 wire _3378_;
 wire _3379_;
 wire _3380_;
 wire _3381_;
 wire _3382_;
 wire _3383_;
 wire _3384_;
 wire _3385_;
 wire _3386_;
 wire _3387_;
 wire _3388_;
 wire _3389_;
 wire _3390_;
 wire _3391_;
 wire _3392_;
 wire _3393_;
 wire _3394_;
 wire _3395_;
 wire _3396_;
 wire _3397_;
 wire _3398_;
 wire _3399_;
 wire _3400_;
 wire _3401_;
 wire _3402_;
 wire _3403_;
 wire _3404_;
 wire _3405_;
 wire _3406_;
 wire _3407_;
 wire _3408_;
 wire _3409_;
 wire _3410_;
 wire _3411_;
 wire _3412_;
 wire _3413_;
 wire _3414_;
 wire _3415_;
 wire _3416_;
 wire _3417_;
 wire _3418_;
 wire _3419_;
 wire _3420_;
 wire _3421_;
 wire _3422_;
 wire _3423_;
 wire _3424_;
 wire _3425_;
 wire _3426_;
 wire _3427_;
 wire _3428_;
 wire _3429_;
 wire _3430_;
 wire _3431_;
 wire _3432_;
 wire _3433_;
 wire _3434_;
 wire _3435_;
 wire _3436_;
 wire _3437_;
 wire _3438_;
 wire _3439_;
 wire _3440_;
 wire _3441_;
 wire _3442_;
 wire _3443_;
 wire _3444_;
 wire _3445_;
 wire _3446_;
 wire _3447_;
 wire _3448_;
 wire _3449_;
 wire _3450_;
 wire _3451_;
 wire _3452_;
 wire _3453_;
 wire _3454_;
 wire _3455_;
 wire _3456_;
 wire _3457_;
 wire _3458_;
 wire _3459_;
 wire _3460_;
 wire _3461_;
 wire _3462_;
 wire _3463_;
 wire _3464_;
 wire _3465_;
 wire _3466_;
 wire _3467_;
 wire _3468_;
 wire _3469_;
 wire _3470_;
 wire _3471_;
 wire _3472_;
 wire _3473_;
 wire _3474_;
 wire _3475_;
 wire _3476_;
 wire _3477_;
 wire _3478_;
 wire _3479_;
 wire _3480_;
 wire _3481_;
 wire _3482_;
 wire _3483_;
 wire _3484_;
 wire _3485_;
 wire _3486_;
 wire _3487_;
 wire _3488_;
 wire _3489_;
 wire _3490_;
 wire _3491_;
 wire _3492_;
 wire _3493_;
 wire _3494_;
 wire _3495_;
 wire _3496_;
 wire _3497_;
 wire _3498_;
 wire _3499_;
 wire _3500_;
 wire _3501_;
 wire _3502_;
 wire _3503_;
 wire _3504_;
 wire _3505_;
 wire _3506_;
 wire _3507_;
 wire _3508_;
 wire _3509_;
 wire _3510_;
 wire _3511_;
 wire _3512_;
 wire _3513_;
 wire _3514_;
 wire _3515_;
 wire _3516_;
 wire _3517_;
 wire _3518_;
 wire _3519_;
 wire _3520_;
 wire _3521_;
 wire _3522_;
 wire _3523_;
 wire _3524_;
 wire _3525_;
 wire _3526_;
 wire _3527_;
 wire _3528_;
 wire _3529_;
 wire _3530_;
 wire _3531_;
 wire _3532_;
 wire _3533_;
 wire _3534_;
 wire _3535_;
 wire _3536_;
 wire _3537_;
 wire _3538_;
 wire _3539_;
 wire _3540_;
 wire _3541_;
 wire _3542_;
 wire _3543_;
 wire _3544_;
 wire _3545_;
 wire _3546_;
 wire _3547_;
 wire _3548_;
 wire _3549_;
 wire _3550_;
 wire _3551_;
 wire _3552_;
 wire _3553_;
 wire _3554_;
 wire _3555_;
 wire _3556_;
 wire _3557_;
 wire _3558_;
 wire _3559_;
 wire _3560_;
 wire _3561_;
 wire _3562_;
 wire _3563_;
 wire _3564_;
 wire _3565_;
 wire _3566_;
 wire _3567_;
 wire _3568_;
 wire _3569_;
 wire _3570_;
 wire _3571_;
 wire _3572_;
 wire _3573_;
 wire _3574_;
 wire _3575_;
 wire _3576_;
 wire _3577_;
 wire _3578_;
 wire _3579_;
 wire _3580_;
 wire _3581_;
 wire _3582_;
 wire _3583_;
 wire _3584_;
 wire _3585_;
 wire _3586_;
 wire _3587_;
 wire _3588_;
 wire _3589_;
 wire _3590_;
 wire _3591_;
 wire _3592_;
 wire _3593_;
 wire _3594_;
 wire _3595_;
 wire _3596_;
 wire _3597_;
 wire _3598_;
 wire _3599_;
 wire _3600_;
 wire _3601_;
 wire _3602_;
 wire _3603_;
 wire _3604_;
 wire _3605_;
 wire _3606_;
 wire _3607_;
 wire _3608_;
 wire _3609_;
 wire _3610_;
 wire _3611_;
 wire _3612_;
 wire _3613_;
 wire _3614_;
 wire _3615_;
 wire _3616_;
 wire _3617_;
 wire _3618_;
 wire _3619_;
 wire _3620_;
 wire _3621_;
 wire _3622_;
 wire _3623_;
 wire _3624_;
 wire _3625_;
 wire _3626_;
 wire _3627_;
 wire _3628_;
 wire _3629_;
 wire _3630_;
 wire _3631_;
 wire _3632_;
 wire _3633_;
 wire _3634_;
 wire _3635_;
 wire _3636_;
 wire _3637_;
 wire _3638_;
 wire _3639_;
 wire _3640_;
 wire _3641_;
 wire _3642_;
 wire _3643_;
 wire _3644_;
 wire _3645_;
 wire _3646_;
 wire _3647_;
 wire _3648_;
 wire _3649_;
 wire _3650_;
 wire _3651_;
 wire _3652_;
 wire _3653_;
 wire _3654_;
 wire _3655_;
 wire _3656_;
 wire _3657_;
 wire _3658_;
 wire _3659_;
 wire _3660_;
 wire _3661_;
 wire _3662_;
 wire _3663_;
 wire _3664_;
 wire _3665_;
 wire _3666_;
 wire _3667_;
 wire _3668_;
 wire _3669_;
 wire _3670_;
 wire _3671_;
 wire _3672_;
 wire _3673_;
 wire _3674_;
 wire _3675_;
 wire _3676_;
 wire _3677_;
 wire _3678_;
 wire _3679_;
 wire _3680_;
 wire _3681_;
 wire _3682_;
 wire _3683_;
 wire _3684_;
 wire _3685_;
 wire _3686_;
 wire _3687_;
 wire _3688_;
 wire _3689_;
 wire _3690_;
 wire _3691_;
 wire _3692_;
 wire _3693_;
 wire _3694_;
 wire _3695_;
 wire _3696_;
 wire _3697_;
 wire _3698_;
 wire _3699_;
 wire _3700_;
 wire _3701_;
 wire _3702_;
 wire _3703_;
 wire _3704_;
 wire _3705_;
 wire _3706_;
 wire _3707_;
 wire _3708_;
 wire _3709_;
 wire _3710_;
 wire _3711_;
 wire _3712_;
 wire _3713_;
 wire _3714_;
 wire _3715_;
 wire _3716_;
 wire _3717_;
 wire _3718_;
 wire _3719_;
 wire _3720_;
 wire _3721_;
 wire _3722_;
 wire _3723_;
 wire _3724_;
 wire _3725_;
 wire _3726_;
 wire _3727_;
 wire _3728_;
 wire _3729_;
 wire _3730_;
 wire _3731_;
 wire _3732_;
 wire _3733_;
 wire _3734_;
 wire _3735_;
 wire _3736_;
 wire _3737_;
 wire _3738_;
 wire _3739_;
 wire _3740_;
 wire _3741_;
 wire _3742_;
 wire _3743_;
 wire _3744_;
 wire _3745_;
 wire _3746_;
 wire _3747_;
 wire _3748_;
 wire _3749_;
 wire _3750_;
 wire _3751_;
 wire _3752_;
 wire _3753_;
 wire _3754_;
 wire _3755_;
 wire _3756_;
 wire _3757_;
 wire _3758_;
 wire _3759_;
 wire _3760_;
 wire _3761_;
 wire _3762_;
 wire _3763_;
 wire _3764_;
 wire _3765_;
 wire _3766_;
 wire _3767_;
 wire _3768_;
 wire _3769_;
 wire _3770_;
 wire _3771_;
 wire _3772_;
 wire _3773_;
 wire _3774_;
 wire _3775_;
 wire _3776_;
 wire _3777_;
 wire _3778_;
 wire _3779_;
 wire _3780_;
 wire _3781_;
 wire _3782_;
 wire _3783_;
 wire _3784_;
 wire _3785_;
 wire _3786_;
 wire _3787_;
 wire _3788_;
 wire _3789_;
 wire _3790_;
 wire _3791_;
 wire _3792_;
 wire _3793_;
 wire _3794_;
 wire _3795_;
 wire _3796_;
 wire _3797_;
 wire _3798_;
 wire _3799_;
 wire _3800_;
 wire _3801_;
 wire _3802_;
 wire _3803_;
 wire _3804_;
 wire _3805_;
 wire _3806_;
 wire _3807_;
 wire _3808_;
 wire _3809_;
 wire _3810_;
 wire _3811_;
 wire _3812_;
 wire _3813_;
 wire _3814_;
 wire _3815_;
 wire _3816_;
 wire _3817_;
 wire _3818_;
 wire _3819_;
 wire _3820_;
 wire _3821_;
 wire _3822_;
 wire _3823_;
 wire _3824_;
 wire _3825_;
 wire _3826_;
 wire _3827_;
 wire _3828_;
 wire _3829_;
 wire _3830_;
 wire _3831_;
 wire _3832_;
 wire _3833_;
 wire _3834_;
 wire _3835_;
 wire _3836_;
 wire _3837_;
 wire _3838_;
 wire _3839_;
 wire _3840_;
 wire _3841_;
 wire _3842_;
 wire _3843_;
 wire _3844_;
 wire _3845_;
 wire _3846_;
 wire _3847_;
 wire _3848_;
 wire _3849_;
 wire _3850_;
 wire _3851_;
 wire _3852_;
 wire _3853_;
 wire _3854_;
 wire _3855_;
 wire _3856_;
 wire _3857_;
 wire _3858_;
 wire _3859_;
 wire _3860_;
 wire _3861_;
 wire _3862_;
 wire _3863_;
 wire _3864_;
 wire _3865_;
 wire _3866_;
 wire _3867_;
 wire _3868_;
 wire _3869_;
 wire _3870_;
 wire _3871_;
 wire _3872_;
 wire _3873_;
 wire _3874_;
 wire _3875_;
 wire _3876_;
 wire _3877_;
 wire _3878_;
 wire _3879_;
 wire _3880_;
 wire _3881_;
 wire _3882_;
 wire _3883_;
 wire _3884_;
 wire _3885_;
 wire _3886_;
 wire _3887_;
 wire _3888_;
 wire _3889_;
 wire _3890_;
 wire _3891_;
 wire _3892_;
 wire _3893_;
 wire _3894_;
 wire _3895_;
 wire _3896_;
 wire _3897_;
 wire _3898_;
 wire _3899_;
 wire _3900_;
 wire _3901_;
 wire _3902_;
 wire _3903_;
 wire _3904_;
 wire _3905_;
 wire _3906_;
 wire _3907_;
 wire _3908_;
 wire _3909_;
 wire _3910_;
 wire _3911_;
 wire _3912_;
 wire _3913_;
 wire _3914_;
 wire _3915_;
 wire _3916_;
 wire _3917_;
 wire _3918_;
 wire _3919_;
 wire _3920_;
 wire _3921_;
 wire _3922_;
 wire _3923_;
 wire _3924_;
 wire _3925_;
 wire _3926_;
 wire _3927_;
 wire _3928_;
 wire _3929_;
 wire _3930_;
 wire _3931_;
 wire _3932_;
 wire _3933_;
 wire _3934_;
 wire _3935_;
 wire _3936_;
 wire _3937_;
 wire _3938_;
 wire _3939_;
 wire _3940_;
 wire _3941_;
 wire _3942_;
 wire _3943_;
 wire _3944_;
 wire _3945_;
 wire _3946_;
 wire _3947_;
 wire _3948_;
 wire _3949_;
 wire _3950_;
 wire _3951_;
 wire _3952_;
 wire _3953_;
 wire _3954_;
 wire _3955_;
 wire _3956_;
 wire _3957_;
 wire _3958_;
 wire _3959_;
 wire _3960_;
 wire _3961_;
 wire _3962_;
 wire _3963_;
 wire _3964_;
 wire _3965_;
 wire _3966_;
 wire _3967_;
 wire _3968_;
 wire _3969_;
 wire _3970_;
 wire _3971_;
 wire _3972_;
 wire _3973_;
 wire _3974_;
 wire _3975_;
 wire _3976_;
 wire _3977_;
 wire _3978_;
 wire _3979_;
 wire _3980_;
 wire _3981_;
 wire _3982_;
 wire _3983_;
 wire _3984_;
 wire _3985_;
 wire _3986_;
 wire _3987_;
 wire _3988_;
 wire _3989_;
 wire _3990_;
 wire _3991_;
 wire _3992_;
 wire _3993_;
 wire _3994_;
 wire _3995_;
 wire _3996_;
 wire _3997_;
 wire _3998_;
 wire _3999_;
 wire _4000_;
 wire _4001_;
 wire _4002_;
 wire _4003_;
 wire _4004_;
 wire _4005_;
 wire _4006_;
 wire _4007_;
 wire _4008_;
 wire _4009_;
 wire _4010_;
 wire _4011_;
 wire _4012_;
 wire _4013_;
 wire _4014_;
 wire _4015_;
 wire _4016_;
 wire _4017_;
 wire _4018_;
 wire _4019_;
 wire _4020_;
 wire _4021_;
 wire _4022_;
 wire _4023_;
 wire _4024_;
 wire _4025_;
 wire _4026_;
 wire _4027_;
 wire _4028_;
 wire _4029_;
 wire _4030_;
 wire _4031_;
 wire _4032_;
 wire _4033_;
 wire _4034_;
 wire _4035_;
 wire _4036_;
 wire _4037_;
 wire _4038_;
 wire _4039_;
 wire _4040_;
 wire _4041_;
 wire _4042_;
 wire _4043_;
 wire _4044_;
 wire _4045_;
 wire _4046_;
 wire _4047_;
 wire _4048_;
 wire _4049_;
 wire _4050_;
 wire _4051_;
 wire _4052_;
 wire _4053_;
 wire _4054_;
 wire _4055_;
 wire _4056_;
 wire _4057_;
 wire _4058_;
 wire _4059_;
 wire _4060_;
 wire _4061_;
 wire _4062_;
 wire _4063_;
 wire _4064_;
 wire _4065_;
 wire _4066_;
 wire _4067_;
 wire _4068_;
 wire _4069_;
 wire _4070_;
 wire _4071_;
 wire _4072_;
 wire _4073_;
 wire _4074_;
 wire _4075_;
 wire _4076_;
 wire _4077_;
 wire _4078_;
 wire _4079_;
 wire _4080_;
 wire _4081_;
 wire _4082_;
 wire _4083_;
 wire _4084_;
 wire _4085_;
 wire _4086_;
 wire _4087_;
 wire _4088_;
 wire _4089_;
 wire _4090_;
 wire _4091_;
 wire _4092_;
 wire _4093_;
 wire _4094_;
 wire _4095_;
 wire _4096_;
 wire _4097_;
 wire _4098_;
 wire _4099_;
 wire _4100_;
 wire _4101_;
 wire _4102_;
 wire _4103_;
 wire _4104_;
 wire _4105_;
 wire _4106_;
 wire _4107_;
 wire _4108_;
 wire _4109_;
 wire _4110_;
 wire _4111_;
 wire _4112_;
 wire _4113_;
 wire _4114_;
 wire _4115_;
 wire _4116_;
 wire _4117_;
 wire _4118_;
 wire _4119_;
 wire _4120_;
 wire _4121_;
 wire _4122_;
 wire _4123_;
 wire _4124_;
 wire _4125_;
 wire _4126_;
 wire _4127_;
 wire _4128_;
 wire _4129_;
 wire _4130_;
 wire _4131_;
 wire _4132_;
 wire _4133_;
 wire _4134_;
 wire _4135_;
 wire _4136_;
 wire _4137_;
 wire _4138_;
 wire _4139_;
 wire _4140_;
 wire _4141_;
 wire _4142_;
 wire _4143_;
 wire _4144_;
 wire _4145_;
 wire _4146_;
 wire _4147_;
 wire _4148_;
 wire _4149_;
 wire _4150_;
 wire _4151_;
 wire _4152_;
 wire _4153_;
 wire _4154_;
 wire _4155_;
 wire _4156_;
 wire _4157_;
 wire _4158_;
 wire _4159_;
 wire _4160_;
 wire _4161_;
 wire _4162_;
 wire _4163_;
 wire _4164_;
 wire _4165_;
 wire _4166_;
 wire _4167_;
 wire _4168_;
 wire _4169_;
 wire _4170_;
 wire _4171_;
 wire _4172_;
 wire _4173_;
 wire _4174_;
 wire _4175_;
 wire _4176_;
 wire _4177_;
 wire _4178_;
 wire _4179_;
 wire _4180_;
 wire _4181_;
 wire _4182_;
 wire _4183_;
 wire _4184_;
 wire _4185_;
 wire _4186_;
 wire _4187_;
 wire _4188_;
 wire _4189_;
 wire _4190_;
 wire _4191_;
 wire _4192_;
 wire _4193_;
 wire _4194_;
 wire _4195_;
 wire _4196_;
 wire _4197_;
 wire _4198_;
 wire _4199_;
 wire _4200_;
 wire _4201_;
 wire _4202_;
 wire _4203_;
 wire _4204_;
 wire _4205_;
 wire _4206_;
 wire _4207_;
 wire _4208_;
 wire _4209_;
 wire _4210_;
 wire _4211_;
 wire _4212_;
 wire _4213_;
 wire _4214_;
 wire _4215_;
 wire _4216_;
 wire _4217_;
 wire _4218_;
 wire _4219_;
 wire _4220_;
 wire _4221_;
 wire _4222_;
 wire _4223_;
 wire _4224_;
 wire _4225_;
 wire _4226_;
 wire _4227_;
 wire _4228_;
 wire _4229_;
 wire _4230_;
 wire _4231_;
 wire _4232_;
 wire _4233_;
 wire _4234_;
 wire _4235_;
 wire _4236_;
 wire _4237_;
 wire _4238_;
 wire _4239_;
 wire _4240_;
 wire _4241_;
 wire _4242_;
 wire _4243_;
 wire _4244_;
 wire _4245_;
 wire _4246_;
 wire _4247_;
 wire _4248_;
 wire _4249_;
 wire _4250_;
 wire _4251_;
 wire _4252_;
 wire _4253_;
 wire _4254_;
 wire _4255_;
 wire _4256_;
 wire _4257_;
 wire _4258_;
 wire _4259_;
 wire _4260_;
 wire _4261_;
 wire _4262_;
 wire _4263_;
 wire _4264_;
 wire _4265_;
 wire _4266_;
 wire _4267_;
 wire _4268_;
 wire _4269_;
 wire _4270_;
 wire _4271_;
 wire _4272_;
 wire _4273_;
 wire _4274_;
 wire _4275_;
 wire _4276_;
 wire _4277_;
 wire _4278_;
 wire _4279_;
 wire _4280_;
 wire _4281_;
 wire _4282_;
 wire _4283_;
 wire _4284_;
 wire _4285_;
 wire _4286_;
 wire _4287_;
 wire _4288_;
 wire _4289_;
 wire _4290_;
 wire _4291_;
 wire _4292_;
 wire _4293_;
 wire _4294_;
 wire _4295_;
 wire _4296_;
 wire _4297_;
 wire _4298_;
 wire _4299_;
 wire _4300_;
 wire _4301_;
 wire _4302_;
 wire _4303_;
 wire _4304_;
 wire _4305_;
 wire _4306_;
 wire _4307_;
 wire _4308_;
 wire _4309_;
 wire _4310_;
 wire _4311_;
 wire _4312_;
 wire _4313_;
 wire _4314_;
 wire _4315_;
 wire _4316_;
 wire _4317_;
 wire _4318_;
 wire _4319_;
 wire _4320_;
 wire _4321_;
 wire _4322_;
 wire _4323_;
 wire _4324_;
 wire _4325_;
 wire _4326_;
 wire _4327_;
 wire _4328_;
 wire _4329_;
 wire _4330_;
 wire _4331_;
 wire _4332_;
 wire _4333_;
 wire _4334_;
 wire _4335_;
 wire _4336_;
 wire _4337_;
 wire _4338_;
 wire _4339_;
 wire _4340_;
 wire _4341_;
 wire _4342_;
 wire _4343_;
 wire _4344_;
 wire _4345_;
 wire _4346_;
 wire _4347_;
 wire _4348_;
 wire _4349_;
 wire _4350_;
 wire _4351_;
 wire _4352_;
 wire _4353_;
 wire _4354_;
 wire _4355_;
 wire _4356_;
 wire _4357_;
 wire _4358_;
 wire _4359_;
 wire _4360_;
 wire _4361_;
 wire _4362_;
 wire _4363_;
 wire _4364_;
 wire _4365_;
 wire _4366_;
 wire _4367_;
 wire _4368_;
 wire _4369_;
 wire _4370_;
 wire _4371_;
 wire _4372_;
 wire _4373_;
 wire _4374_;
 wire _4375_;
 wire _4376_;
 wire _4377_;
 wire _4378_;
 wire _4379_;
 wire _4380_;
 wire _4381_;
 wire _4382_;
 wire _4383_;
 wire _4384_;
 wire _4385_;
 wire _4386_;
 wire _4387_;
 wire _4388_;
 wire _4389_;
 wire _4390_;
 wire _4391_;
 wire _4392_;
 wire _4393_;
 wire _4394_;
 wire _4395_;
 wire _4396_;
 wire _4397_;
 wire _4398_;
 wire _4399_;
 wire _4400_;
 wire _4401_;
 wire _4402_;
 wire _4403_;
 wire _4404_;
 wire _4405_;
 wire _4406_;
 wire _4407_;
 wire _4408_;
 wire _4409_;
 wire _4410_;
 wire _4411_;
 wire _4412_;
 wire _4413_;
 wire _4414_;
 wire _4415_;
 wire _4416_;
 wire _4417_;
 wire _4418_;
 wire _4419_;
 wire _4420_;
 wire _4421_;
 wire _4422_;
 wire _4423_;
 wire _4424_;
 wire _4425_;
 wire _4426_;
 wire _4427_;
 wire _4428_;
 wire _4429_;
 wire _4430_;
 wire _4431_;
 wire _4432_;
 wire _4433_;
 wire _4434_;
 wire _4435_;
 wire _4436_;
 wire _4437_;
 wire _4438_;
 wire _4439_;
 wire _4440_;
 wire _4441_;
 wire _4442_;
 wire _4443_;
 wire _4444_;
 wire _4445_;
 wire _4446_;
 wire _4447_;
 wire _4448_;
 wire _4449_;
 wire _4450_;
 wire _4451_;
 wire _4452_;
 wire _4453_;
 wire _4454_;
 wire _4455_;
 wire _4456_;
 wire _4457_;
 wire _4458_;
 wire _4459_;
 wire _4460_;
 wire _4461_;
 wire _4462_;
 wire _4463_;
 wire _4464_;
 wire _4465_;
 wire _4466_;
 wire _4467_;
 wire _4468_;
 wire _4469_;
 wire _4470_;
 wire _4471_;
 wire _4472_;
 wire _4473_;
 wire _4474_;
 wire _4475_;
 wire _4476_;
 wire _4477_;
 wire _4478_;
 wire _4479_;
 wire _4480_;
 wire _4481_;
 wire _4482_;
 wire _4483_;
 wire _4484_;
 wire _4485_;
 wire _4486_;
 wire _4487_;
 wire _4488_;
 wire _4489_;
 wire _4490_;
 wire _4491_;
 wire _4492_;
 wire _4493_;
 wire _4494_;
 wire _4495_;
 wire _4496_;
 wire _4497_;
 wire _4498_;
 wire _4499_;
 wire _4500_;
 wire _4501_;
 wire _4502_;
 wire _4503_;
 wire _4504_;
 wire _4505_;
 wire _4506_;
 wire _4507_;
 wire _4508_;
 wire _4509_;
 wire _4510_;
 wire _4511_;
 wire _4512_;
 wire _4513_;
 wire _4514_;
 wire _4515_;
 wire _4516_;
 wire _4517_;
 wire _4518_;
 wire _4519_;
 wire _4520_;
 wire _4521_;
 wire _4522_;
 wire _4523_;
 wire _4524_;
 wire _4525_;
 wire _4526_;
 wire _4527_;
 wire _4528_;
 wire _4529_;
 wire _4530_;
 wire _4531_;
 wire _4532_;
 wire _4533_;
 wire _4534_;
 wire _4535_;
 wire _4536_;
 wire _4537_;
 wire _4538_;
 wire _4539_;
 wire _4540_;
 wire _4541_;
 wire _4542_;
 wire _4543_;
 wire _4544_;
 wire _4545_;
 wire _4546_;
 wire _4547_;
 wire _4548_;
 wire _4549_;
 wire _4550_;
 wire _4551_;
 wire _4552_;
 wire \as2650.addr_buff[0] ;
 wire \as2650.addr_buff[1] ;
 wire \as2650.addr_buff[2] ;
 wire \as2650.addr_buff[3] ;
 wire \as2650.addr_buff[4] ;
 wire \as2650.addr_buff[5] ;
 wire \as2650.addr_buff[6] ;
 wire \as2650.addr_buff[7] ;
 wire \as2650.carry ;
 wire \as2650.cycle[0] ;
 wire \as2650.cycle[1] ;
 wire \as2650.cycle[2] ;
 wire \as2650.cycle[3] ;
 wire \as2650.cycle[4] ;
 wire \as2650.cycle[5] ;
 wire \as2650.cycle[6] ;
 wire \as2650.cycle[7] ;
 wire \as2650.halted ;
 wire \as2650.holding_reg[0] ;
 wire \as2650.holding_reg[1] ;
 wire \as2650.holding_reg[2] ;
 wire \as2650.holding_reg[3] ;
 wire \as2650.holding_reg[4] ;
 wire \as2650.holding_reg[5] ;
 wire \as2650.holding_reg[6] ;
 wire \as2650.holding_reg[7] ;
 wire \as2650.idx_ctrl[0] ;
 wire \as2650.idx_ctrl[1] ;
 wire \as2650.ins_reg[0] ;
 wire \as2650.ins_reg[1] ;
 wire \as2650.ins_reg[2] ;
 wire \as2650.ins_reg[3] ;
 wire \as2650.ins_reg[4] ;
 wire \as2650.ins_reg[5] ;
 wire \as2650.ins_reg[6] ;
 wire \as2650.ins_reg[7] ;
 wire \as2650.overflow ;
 wire \as2650.pc[0] ;
 wire \as2650.pc[10] ;
 wire \as2650.pc[11] ;
 wire \as2650.pc[12] ;
 wire \as2650.pc[13] ;
 wire \as2650.pc[14] ;
 wire \as2650.pc[1] ;
 wire \as2650.pc[2] ;
 wire \as2650.pc[3] ;
 wire \as2650.pc[4] ;
 wire \as2650.pc[5] ;
 wire \as2650.pc[6] ;
 wire \as2650.pc[7] ;
 wire \as2650.pc[8] ;
 wire \as2650.pc[9] ;
 wire \as2650.psl[1] ;
 wire \as2650.psl[3] ;
 wire \as2650.psl[4] ;
 wire \as2650.psl[5] ;
 wire \as2650.psl[6] ;
 wire \as2650.psl[7] ;
 wire \as2650.psu[0] ;
 wire \as2650.psu[1] ;
 wire \as2650.psu[2] ;
 wire \as2650.psu[3] ;
 wire \as2650.psu[4] ;
 wire \as2650.psu[5] ;
 wire \as2650.psu[7] ;
 wire \as2650.r0[0] ;
 wire \as2650.r0[1] ;
 wire \as2650.r0[2] ;
 wire \as2650.r0[3] ;
 wire \as2650.r0[4] ;
 wire \as2650.r0[5] ;
 wire \as2650.r0[6] ;
 wire \as2650.r0[7] ;
 wire \as2650.r123[0][0] ;
 wire \as2650.r123[0][1] ;
 wire \as2650.r123[0][2] ;
 wire \as2650.r123[0][3] ;
 wire \as2650.r123[0][4] ;
 wire \as2650.r123[0][5] ;
 wire \as2650.r123[0][6] ;
 wire \as2650.r123[0][7] ;
 wire \as2650.r123[1][0] ;
 wire \as2650.r123[1][1] ;
 wire \as2650.r123[1][2] ;
 wire \as2650.r123[1][3] ;
 wire \as2650.r123[1][4] ;
 wire \as2650.r123[1][5] ;
 wire \as2650.r123[1][6] ;
 wire \as2650.r123[1][7] ;
 wire \as2650.r123[2][0] ;
 wire \as2650.r123[2][1] ;
 wire \as2650.r123[2][2] ;
 wire \as2650.r123[2][3] ;
 wire \as2650.r123[2][4] ;
 wire \as2650.r123[2][5] ;
 wire \as2650.r123[2][6] ;
 wire \as2650.r123[2][7] ;
 wire \as2650.r123[3][0] ;
 wire \as2650.r123[3][1] ;
 wire \as2650.r123[3][2] ;
 wire \as2650.r123[3][3] ;
 wire \as2650.r123[3][4] ;
 wire \as2650.r123[3][5] ;
 wire \as2650.r123[3][6] ;
 wire \as2650.r123[3][7] ;
 wire \as2650.r123_2[0][0] ;
 wire \as2650.r123_2[0][1] ;
 wire \as2650.r123_2[0][2] ;
 wire \as2650.r123_2[0][3] ;
 wire \as2650.r123_2[0][4] ;
 wire \as2650.r123_2[0][5] ;
 wire \as2650.r123_2[0][6] ;
 wire \as2650.r123_2[0][7] ;
 wire \as2650.r123_2[1][0] ;
 wire \as2650.r123_2[1][1] ;
 wire \as2650.r123_2[1][2] ;
 wire \as2650.r123_2[1][3] ;
 wire \as2650.r123_2[1][4] ;
 wire \as2650.r123_2[1][5] ;
 wire \as2650.r123_2[1][6] ;
 wire \as2650.r123_2[1][7] ;
 wire \as2650.r123_2[2][0] ;
 wire \as2650.r123_2[2][1] ;
 wire \as2650.r123_2[2][2] ;
 wire \as2650.r123_2[2][3] ;
 wire \as2650.r123_2[2][4] ;
 wire \as2650.r123_2[2][5] ;
 wire \as2650.r123_2[2][6] ;
 wire \as2650.r123_2[2][7] ;
 wire \as2650.r123_2[3][0] ;
 wire \as2650.r123_2[3][1] ;
 wire \as2650.r123_2[3][2] ;
 wire \as2650.r123_2[3][3] ;
 wire \as2650.r123_2[3][4] ;
 wire \as2650.r123_2[3][5] ;
 wire \as2650.r123_2[3][6] ;
 wire \as2650.r123_2[3][7] ;
 wire \as2650.stack[0][0] ;
 wire \as2650.stack[0][10] ;
 wire \as2650.stack[0][11] ;
 wire \as2650.stack[0][12] ;
 wire \as2650.stack[0][13] ;
 wire \as2650.stack[0][14] ;
 wire \as2650.stack[0][1] ;
 wire \as2650.stack[0][2] ;
 wire \as2650.stack[0][3] ;
 wire \as2650.stack[0][4] ;
 wire \as2650.stack[0][5] ;
 wire \as2650.stack[0][6] ;
 wire \as2650.stack[0][7] ;
 wire \as2650.stack[0][8] ;
 wire \as2650.stack[0][9] ;
 wire \as2650.stack[1][0] ;
 wire \as2650.stack[1][10] ;
 wire \as2650.stack[1][11] ;
 wire \as2650.stack[1][12] ;
 wire \as2650.stack[1][13] ;
 wire \as2650.stack[1][14] ;
 wire \as2650.stack[1][1] ;
 wire \as2650.stack[1][2] ;
 wire \as2650.stack[1][3] ;
 wire \as2650.stack[1][4] ;
 wire \as2650.stack[1][5] ;
 wire \as2650.stack[1][6] ;
 wire \as2650.stack[1][7] ;
 wire \as2650.stack[1][8] ;
 wire \as2650.stack[1][9] ;
 wire \as2650.stack[2][0] ;
 wire \as2650.stack[2][10] ;
 wire \as2650.stack[2][11] ;
 wire \as2650.stack[2][12] ;
 wire \as2650.stack[2][13] ;
 wire \as2650.stack[2][14] ;
 wire \as2650.stack[2][1] ;
 wire \as2650.stack[2][2] ;
 wire \as2650.stack[2][3] ;
 wire \as2650.stack[2][4] ;
 wire \as2650.stack[2][5] ;
 wire \as2650.stack[2][6] ;
 wire \as2650.stack[2][7] ;
 wire \as2650.stack[2][8] ;
 wire \as2650.stack[2][9] ;
 wire \as2650.stack[3][0] ;
 wire \as2650.stack[3][10] ;
 wire \as2650.stack[3][11] ;
 wire \as2650.stack[3][12] ;
 wire \as2650.stack[3][13] ;
 wire \as2650.stack[3][14] ;
 wire \as2650.stack[3][1] ;
 wire \as2650.stack[3][2] ;
 wire \as2650.stack[3][3] ;
 wire \as2650.stack[3][4] ;
 wire \as2650.stack[3][5] ;
 wire \as2650.stack[3][6] ;
 wire \as2650.stack[3][7] ;
 wire \as2650.stack[3][8] ;
 wire \as2650.stack[3][9] ;
 wire \as2650.stack[4][0] ;
 wire \as2650.stack[4][10] ;
 wire \as2650.stack[4][11] ;
 wire \as2650.stack[4][12] ;
 wire \as2650.stack[4][13] ;
 wire \as2650.stack[4][14] ;
 wire \as2650.stack[4][1] ;
 wire \as2650.stack[4][2] ;
 wire \as2650.stack[4][3] ;
 wire \as2650.stack[4][4] ;
 wire \as2650.stack[4][5] ;
 wire \as2650.stack[4][6] ;
 wire \as2650.stack[4][7] ;
 wire \as2650.stack[4][8] ;
 wire \as2650.stack[4][9] ;
 wire \as2650.stack[5][0] ;
 wire \as2650.stack[5][10] ;
 wire \as2650.stack[5][11] ;
 wire \as2650.stack[5][12] ;
 wire \as2650.stack[5][13] ;
 wire \as2650.stack[5][14] ;
 wire \as2650.stack[5][1] ;
 wire \as2650.stack[5][2] ;
 wire \as2650.stack[5][3] ;
 wire \as2650.stack[5][4] ;
 wire \as2650.stack[5][5] ;
 wire \as2650.stack[5][6] ;
 wire \as2650.stack[5][7] ;
 wire \as2650.stack[5][8] ;
 wire \as2650.stack[5][9] ;
 wire \as2650.stack[6][0] ;
 wire \as2650.stack[6][10] ;
 wire \as2650.stack[6][11] ;
 wire \as2650.stack[6][12] ;
 wire \as2650.stack[6][13] ;
 wire \as2650.stack[6][14] ;
 wire \as2650.stack[6][1] ;
 wire \as2650.stack[6][2] ;
 wire \as2650.stack[6][3] ;
 wire \as2650.stack[6][4] ;
 wire \as2650.stack[6][5] ;
 wire \as2650.stack[6][6] ;
 wire \as2650.stack[6][7] ;
 wire \as2650.stack[6][8] ;
 wire \as2650.stack[6][9] ;
 wire \as2650.stack[7][0] ;
 wire \as2650.stack[7][10] ;
 wire \as2650.stack[7][11] ;
 wire \as2650.stack[7][12] ;
 wire \as2650.stack[7][13] ;
 wire \as2650.stack[7][14] ;
 wire \as2650.stack[7][1] ;
 wire \as2650.stack[7][2] ;
 wire \as2650.stack[7][3] ;
 wire \as2650.stack[7][4] ;
 wire \as2650.stack[7][5] ;
 wire \as2650.stack[7][6] ;
 wire \as2650.stack[7][7] ;
 wire \as2650.stack[7][8] ;
 wire \as2650.stack[7][9] ;
 wire clknet_0_wb_clk_i;
 wire clknet_3_0_0_wb_clk_i;
 wire clknet_3_1_0_wb_clk_i;
 wire clknet_3_2_0_wb_clk_i;
 wire clknet_3_3_0_wb_clk_i;
 wire clknet_3_4_0_wb_clk_i;
 wire clknet_3_5_0_wb_clk_i;
 wire clknet_3_6_0_wb_clk_i;
 wire clknet_3_7_0_wb_clk_i;
 wire clknet_leaf_11_wb_clk_i;
 wire clknet_leaf_12_wb_clk_i;
 wire clknet_leaf_14_wb_clk_i;
 wire clknet_leaf_15_wb_clk_i;
 wire clknet_leaf_16_wb_clk_i;
 wire clknet_leaf_18_wb_clk_i;
 wire clknet_leaf_1_wb_clk_i;
 wire clknet_leaf_20_wb_clk_i;
 wire clknet_leaf_23_wb_clk_i;
 wire clknet_leaf_24_wb_clk_i;
 wire clknet_leaf_25_wb_clk_i;
 wire clknet_leaf_26_wb_clk_i;
 wire clknet_leaf_27_wb_clk_i;
 wire clknet_leaf_28_wb_clk_i;
 wire clknet_leaf_29_wb_clk_i;
 wire clknet_leaf_2_wb_clk_i;
 wire clknet_leaf_30_wb_clk_i;
 wire clknet_leaf_31_wb_clk_i;
 wire clknet_leaf_36_wb_clk_i;
 wire clknet_leaf_37_wb_clk_i;
 wire clknet_leaf_38_wb_clk_i;
 wire clknet_leaf_39_wb_clk_i;
 wire clknet_leaf_3_wb_clk_i;
 wire clknet_leaf_40_wb_clk_i;
 wire clknet_leaf_41_wb_clk_i;
 wire clknet_leaf_42_wb_clk_i;
 wire clknet_leaf_44_wb_clk_i;
 wire clknet_leaf_45_wb_clk_i;
 wire clknet_leaf_46_wb_clk_i;
 wire clknet_leaf_47_wb_clk_i;
 wire clknet_leaf_48_wb_clk_i;
 wire clknet_leaf_49_wb_clk_i;
 wire clknet_leaf_50_wb_clk_i;
 wire clknet_leaf_51_wb_clk_i;
 wire clknet_leaf_52_wb_clk_i;
 wire clknet_leaf_53_wb_clk_i;
 wire clknet_leaf_54_wb_clk_i;
 wire clknet_leaf_55_wb_clk_i;
 wire clknet_leaf_56_wb_clk_i;
 wire clknet_leaf_57_wb_clk_i;
 wire clknet_leaf_58_wb_clk_i;
 wire clknet_leaf_59_wb_clk_i;
 wire clknet_leaf_5_wb_clk_i;
 wire clknet_leaf_60_wb_clk_i;
 wire clknet_leaf_61_wb_clk_i;
 wire clknet_leaf_62_wb_clk_i;
 wire clknet_leaf_63_wb_clk_i;
 wire clknet_leaf_64_wb_clk_i;
 wire clknet_leaf_65_wb_clk_i;
 wire clknet_leaf_66_wb_clk_i;
 wire clknet_leaf_67_wb_clk_i;
 wire clknet_leaf_68_wb_clk_i;
 wire clknet_leaf_69_wb_clk_i;
 wire clknet_leaf_6_wb_clk_i;
 wire clknet_leaf_71_wb_clk_i;
 wire clknet_leaf_73_wb_clk_i;
 wire clknet_leaf_74_wb_clk_i;
 wire clknet_leaf_75_wb_clk_i;
 wire clknet_leaf_76_wb_clk_i;
 wire clknet_leaf_77_wb_clk_i;
 wire clknet_leaf_80_wb_clk_i;
 wire clknet_leaf_8_wb_clk_i;
 wire clknet_leaf_9_wb_clk_i;
 wire clknet_opt_1_0_wb_clk_i;
 wire net1;
 wire net10;
 wire net11;
 wire net12;
 wire net13;
 wire net14;
 wire net15;
 wire net16;
 wire net17;
 wire net18;
 wire net19;
 wire net2;
 wire net20;
 wire net21;
 wire net22;
 wire net23;
 wire net24;
 wire net25;
 wire net26;
 wire net27;
 wire net28;
 wire net29;
 wire net3;
 wire net30;
 wire net31;
 wire net32;
 wire net33;
 wire net34;
 wire net35;
 wire net36;
 wire net37;
 wire net38;
 wire net39;
 wire net4;
 wire net40;
 wire net41;
 wire net42;
 wire net43;
 wire net44;
 wire net45;
 wire net46;
 wire net47;
 wire net48;
 wire net49;
 wire net5;
 wire net50;
 wire net51;
 wire net52;
 wire net53;
 wire net54;
 wire net6;
 wire net7;
 wire net8;
 wire net9;

 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4553__I (.I(net26));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4555__I (.I(_4135_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4557__I (.I(\as2650.ins_reg[0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4558__I (.I(_4138_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4559__A1 (.I(_4139_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4559__A2 (.I(_4135_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4560__I (.I(_4140_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4562__I (.I(_4142_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4564__I (.I(_4144_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4567__I (.I(_4147_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4568__I (.I(_4148_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4570__A2 (.I(net5));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4571__I (.I(_4151_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4572__A2 (.I(_4152_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4573__A1 (.I(_4143_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4573__A2 (.I(_4153_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4575__I (.I(_4155_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4579__I (.I(_4159_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4580__A1 (.I(_4157_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4580__A2 (.I(_4160_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4581__I (.I(\as2650.ins_reg[3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4584__A1 (.I(\as2650.cycle[3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4585__I (.I(_4165_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4586__A1 (.I(_4163_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4587__I (.I(\as2650.cycle[0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4588__A1 (.I(\as2650.cycle[1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4589__A1 (.I(_4167_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4590__A2 (.I(_4170_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4591__I (.I(_4163_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4592__I (.I(\as2650.cycle[1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4594__A1 (.I(_4174_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4595__A1 (.I(_4172_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4595__A3 (.I(_4175_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4600__I (.I(_4180_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4601__I (.I(\as2650.ins_reg[5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4603__A1 (.I(_4155_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4603__A2 (.I(_4183_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4604__A1 (.I(_4181_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4604__A2 (.I(_4184_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4605__A1 (.I(_4179_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4606__A1 (.I(\as2650.ins_reg[3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4607__A1 (.I(_4176_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4607__A2 (.I(_4187_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4608__A1 (.I(_4161_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4608__A2 (.I(_4171_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4608__B (.I(_4188_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4609__A2 (.I(\as2650.ins_reg[3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4610__I (.I(_4190_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4611__I (.I(_4183_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4613__A2 (.I(_4192_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4613__A3 (.I(_4193_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4614__A1 (.I(_4191_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4614__A2 (.I(_4194_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4615__I (.I(_4138_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4616__I (.I(_4196_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4617__A1 (.I(_4197_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4617__A2 (.I(_4135_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4618__I (.I(_4198_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4620__I (.I(_4200_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4621__I (.I(net5));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4622__I (.I(_4202_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4623__A1 (.I(_4201_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4624__A2 (.I(_4204_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4625__A1 (.I(_4199_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4626__A1 (.I(_4163_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4626__A2 (.I(_4165_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4627__I (.I(\as2650.cycle[0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4628__A2 (.I(_4208_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4630__I (.I(_4210_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4631__A1 (.I(_4206_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4631__A2 (.I(_4211_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4632__A1 (.I(_4195_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4632__A2 (.I(_4212_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4634__I (.I(_4181_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4638__A1 (.I(_4215_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4638__A2 (.I(_4218_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4639__A1 (.I(_4214_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4639__A2 (.I(_4219_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4640__A1 (.I(_4212_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4640__A2 (.I(_4220_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4641__I (.I(_4221_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4644__A1 (.I(_4159_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4644__A2 (.I(_4179_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4645__A1 (.I(_4192_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4645__A2 (.I(_4225_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4646__A1 (.I(_4181_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4646__A3 (.I(_4226_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4647__A1 (.I(_4223_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4647__A2 (.I(_4227_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4648__A1 (.I(_4212_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4648__A2 (.I(_4228_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4649__I (.I(_4229_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4652__I (.I(_4232_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4655__A2 (.I(\as2650.cycle[0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4659__A1 (.I(_4238_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4659__A3 (.I(_4165_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4660__A1 (.I(_4237_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4660__A2 (.I(_4240_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4661__A1 (.I(_4235_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4661__A2 (.I(_4241_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4665__I (.I(_4245_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4666__A1 (.I(_4233_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4666__A2 (.I(_4206_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4666__A3 (.I(_4242_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4666__A4 (.I(_4246_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4669__I (.I(_4249_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4670__I (.I(\as2650.cycle[3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4671__A1 (.I(\as2650.cycle[1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4671__A2 (.I(\as2650.cycle[0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4673__A1 (.I(_4163_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4673__A2 (.I(_4253_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4674__I (.I(\as2650.ins_reg[3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4675__A1 (.I(_4181_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4675__A2 (.I(_4255_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4676__I (.I(_4256_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4677__A1 (.I(\as2650.ins_reg[5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4678__A1 (.I(_4198_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4678__A2 (.I(_4257_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4678__A3 (.I(_4245_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4678__A4 (.I(_4258_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4679__A1 (.I(_4254_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4679__A2 (.I(_4259_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4680__A1 (.I(_4250_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4680__A2 (.I(_4151_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4680__A3 (.I(_4260_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4681__A1 (.I(_4248_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4681__A2 (.I(_4261_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4682__A1 (.I(_4235_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4682__A3 (.I(_4240_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4685__A1 (.I(_4264_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4685__A2 (.I(_4265_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4686__A1 (.I(\as2650.addr_buff[7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4687__A1 (.I(_4263_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4688__A1 (.I(_4233_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4688__A2 (.I(_4206_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4688__A3 (.I(_4268_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4689__A1 (.I(_4247_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4689__A2 (.I(_4262_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4689__A3 (.I(_4269_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4690__A1 (.I(_4213_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4690__A3 (.I(_4231_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4691__A1 (.I(_4154_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4691__A2 (.I(_4189_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4691__B (.I(_4271_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4692__A2 (.I(_4272_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4694__I (.I(_4274_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4695__I (.I(_4262_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4696__I (.I(_4192_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4697__A1 (.I(_4159_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4698__A1 (.I(_4277_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4698__A2 (.I(_4278_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4699__A1 (.I(_4138_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4700__S (.I(_4147_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4701__A1 (.I(_4280_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4701__A2 (.I(_4281_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4702__I (.I(_4282_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4703__I (.I(\as2650.r0[0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4704__I (.I(_4284_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4705__A1 (.I(_4138_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4705__A2 (.I(_4135_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4706__I0 (.I(\as2650.r123[1][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4706__I1 (.I(\as2650.r123[0][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4706__I3 (.I(\as2650.r123_2[0][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4706__S0 (.I(\as2650.ins_reg[0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4707__A1 (.I(_4285_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4707__A2 (.I(_4140_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4707__B1 (.I(_4286_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4707__B2 (.I(_4287_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4708__I (.I(_4288_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4709__A1 (.I(_4190_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4711__A1 (.I(_4291_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4711__A2 (.I(_4190_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4713__I (.I(_4285_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4715__A1 (.I(_4295_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4715__A2 (.I(_4198_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4716__I (.I(_4280_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4718__A2 (.I(_4281_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4719__I (.I(_4286_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4720__A2 (.I(_4287_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4721__A1 (.I(_4296_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4721__A2 (.I(_4299_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4721__A3 (.I(_4301_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4721__B (.I(_4291_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4722__A3 (.I(_4302_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4727__A1 (.I(_4305_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4727__A2 (.I(_4306_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4728__A1 (.I(_4291_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4728__A2 (.I(_4256_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4729__A1 (.I(_4256_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4729__A2 (.I(_4304_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4730__A1 (.I(_4303_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4730__A2 (.I(_4310_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4731__I (.I(_4183_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4732__A1 (.I(_4159_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4732__A2 (.I(_4179_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4733__I (.I(_4313_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4734__A1 (.I(_4312_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4734__A2 (.I(_4314_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4735__I (.I(\as2650.carry ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4736__A1 (.I(\as2650.psl[3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4736__A2 (.I(_4316_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4737__A2 (.I(_4311_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4738__A1 (.I(_4315_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4739__I (.I(\as2650.psl[3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4740__A1 (.I(_4320_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4740__A2 (.I(\as2650.carry ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4741__A1 (.I(_4321_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4741__A2 (.I(_4311_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4742__I (.I(_4160_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4743__A1 (.I(_4323_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4744__A1 (.I(_4192_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4744__A2 (.I(_4324_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4745__A1 (.I(_4303_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4745__A2 (.I(_4310_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4745__B (.I(\as2650.psl[3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4745__C (.I(\as2650.carry ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4746__A2 (.I(_4325_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4748__A1 (.I(_4323_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4748__A2 (.I(_4328_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4749__I (.I(_4329_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4750__I (.I(_4257_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4752__I (.I(_4304_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4753__I (.I(_4333_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4754__A1 (.I(_4332_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4754__A2 (.I(_4334_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4755__I (.I(_4324_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4757__I (.I(_4226_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4758__A1 (.I(_4330_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4758__B1 (.I(_4336_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4758__C (.I(_4338_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4760__A1 (.I(_4183_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4760__A2 (.I(_4225_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4761__A1 (.I(_4341_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4761__B (.I(_4279_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4762__A1 (.I(_4279_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4762__A2 (.I(_4311_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4764__I (.I(_4247_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4765__I (.I(_4345_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4770__A1 (.I(_4348_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4770__A2 (.I(_4350_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4771__A1 (.I(_4304_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4772__I (.I(_4352_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4773__I (.I(_4269_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4777__A1 (.I(_4357_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4779__A1 (.I(_4333_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4779__A2 (.I(_4359_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4781__I (.I(_4213_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4783__I (.I(_4221_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4784__I (.I(_4320_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4787__A1 (.I(_4367_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4787__A2 (.I(_4142_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4789__S (.I(_4148_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4790__A1 (.I(_4369_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4790__A2 (.I(_4370_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4791__I1 (.I(\as2650.r123[0][7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4791__I3 (.I(\as2650.r123_2[0][7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4791__S0 (.I(_4197_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4791__S1 (.I(_4148_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4792__A2 (.I(_4372_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4793__A1 (.I(_4368_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4794__I (.I(_4374_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4795__I (.I(_4375_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4796__A1 (.I(_4365_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4796__A2 (.I(_4376_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4796__B (.I(_4321_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4799__S (.I(_4379_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4800__A2 (.I(_4380_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4802__I (.I(_4382_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4803__I1 (.I(\as2650.r123[0][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4803__I2 (.I(\as2650.r123_2[1][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4803__I3 (.I(\as2650.r123_2[0][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4803__S0 (.I(_4139_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4803__S1 (.I(_4379_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4804__A1 (.I(_4383_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4804__A2 (.I(_4140_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4804__B1 (.I(_4286_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4804__B2 (.I(_4384_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4805__A1 (.I(_4381_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4805__A2 (.I(_4385_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4806__I (.I(_4386_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4807__I (.I(_4387_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4808__I (.I(_4229_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4809__I (.I(net6));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4810__I (.I(_4390_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4811__I (.I(_4391_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4812__A1 (.I(_4172_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4812__A3 (.I(_4175_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4814__A2 (.I(_4393_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4814__A3 (.I(_4394_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4815__A1 (.I(_4154_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4815__A2 (.I(_4395_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4816__I (.I(_4396_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4817__A2 (.I(_4333_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4818__I (.I(_4396_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4819__A1 (.I(_4398_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4819__A2 (.I(_4399_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4820__A1 (.I(_4392_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4822__A1 (.I(_4378_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4822__A2 (.I(_4388_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4823__A2 (.I(_4377_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4823__B (.I(_4403_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4824__I (.I(_4285_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4825__I (.I(_4405_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4826__A1 (.I(_4157_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4826__A2 (.I(_4268_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4827__A1 (.I(_4154_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4828__A1 (.I(_4406_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4828__B (.I(_4408_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4830__A1 (.I(_4354_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4830__A2 (.I(_4361_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4830__C (.I(_4345_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4831__I (.I(_4262_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4832__A2 (.I(_4353_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4833__A2 (.I(_4344_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4835__I (.I(_4415_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4836__I (.I(_4170_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4837__I (.I(_4417_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4838__I (.I(_4418_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4839__I (.I(_4143_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4840__I (.I(_4190_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4842__A2 (.I(_4278_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4843__A1 (.I(_4312_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4843__A2 (.I(_4423_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4845__A1 (.I(_4420_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4845__A2 (.I(_4422_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4845__A3 (.I(_4425_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4847__I (.I(_4197_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4848__A1 (.I(_4428_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4850__A2 (.I(_4313_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4851__A1 (.I(_4312_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4851__A2 (.I(_4431_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4852__A1 (.I(_4427_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4852__A2 (.I(_4430_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4852__A3 (.I(_4432_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4853__A1 (.I(_4426_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4854__I (.I(_4434_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4855__A1 (.I(_4419_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4855__A2 (.I(_4435_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4857__I (.I(_4202_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4858__C (.I(_4438_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4860__I (.I(_4406_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4861__I (.I(_4211_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4862__I (.I(_4442_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4863__A1 (.I(_4443_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4863__A2 (.I(_4426_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4864__A1 (.I(_4415_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4864__A2 (.I(_4444_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4865__I (.I(_4445_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4866__A1 (.I(_4441_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4870__A2 (.I(_4450_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4873__I (.I(_4453_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4874__A2 (.I(_4452_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4874__B (.I(_4454_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4878__A2 (.I(_4458_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4880__I (.I(_4460_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4881__A1 (.I(\as2650.stack[2][8] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4881__A2 (.I(_4461_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4883__A2 (.I(_4463_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4885__I (.I(_4465_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4887__A2 (.I(_4458_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4889__I (.I(_4469_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4890__A2 (.I(_4466_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4890__B1 (.I(_4470_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4891__A2 (.I(_4462_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4892__A2 (.I(_4450_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4894__A1 (.I(_4473_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4894__A2 (.I(_4474_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4895__I (.I(_4475_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4896__I (.I(_4476_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4897__I (.I(_4450_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4898__I (.I(_4478_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4899__A2 (.I(_4479_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4899__B1 (.I(_4461_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4901__I (.I(_4481_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4902__A2 (.I(_4482_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4902__B1 (.I(_4470_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4903__A1 (.I(_4477_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4904__I (.I(_4445_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4905__A1 (.I(_4472_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4905__A2 (.I(_4484_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4906__I (.I(_4211_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4907__I (.I(_4191_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4908__A1 (.I(_4143_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4908__A2 (.I(_4488_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4908__A3 (.I(_4432_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4909__A2 (.I(_4489_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4910__I (.I(_4490_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4911__A2 (.I(_4491_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4912__A1 (.I(_4415_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4914__A3 (.I(_4486_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4914__A4 (.I(_4494_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4915__A1 (.I(\as2650.r123[0][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4916__A2 (.I(_4414_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4917__I (.I(\as2650.r123[0][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4920__I (.I(_4274_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4921__I (.I(_4408_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4924__A1 (.I(_4305_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4924__A2 (.I(_4306_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4924__A3 (.I(_4503_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4925__B1 (.I(_4381_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4925__B2 (.I(_4385_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4926__I (.I(_4505_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4927__I (.I(_4506_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4928__A1 (.I(_4282_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4928__A2 (.I(_4288_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4928__A3 (.I(_4381_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4928__A4 (.I(_4385_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4929__I (.I(_4508_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4930__I (.I(_4509_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4931__A3 (.I(_4507_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4931__A4 (.I(_4510_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4932__B1 (.I(_4507_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4932__B2 (.I(_4510_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4933__A1 (.I(_4511_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4933__A2 (.I(_4512_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4934__A1 (.I(_4305_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4934__A2 (.I(_4306_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4936__I (.I(_4147_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4937__S (.I(_4516_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4938__A2 (.I(_4517_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4939__I (.I(\as2650.r0[2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4940__I (.I(_4519_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4941__I (.I(_4286_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4942__I1 (.I(\as2650.r123[0][2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4942__I3 (.I(\as2650.r123_2[0][2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4942__S0 (.I(_4139_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4942__S1 (.I(_4379_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4943__A1 (.I(_4520_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4943__A2 (.I(_4140_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4943__B1 (.I(_4521_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4943__B2 (.I(_4522_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4944__A1 (.I(_4518_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4944__A2 (.I(_4523_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4945__I (.I(_4524_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4946__I (.I(_4525_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4947__I (.I(_4526_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4948__I (.I(net7));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4949__I (.I(_4528_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4950__I (.I(_4529_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4951__I (.I(_4530_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4952__I (.I(_4399_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4953__A1 (.I(_4249_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4953__A2 (.I(_4258_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4954__I1 (.I(_4533_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4954__S (.I(_4333_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4955__A1 (.I(_4387_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4955__A2 (.I(_4534_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4956__A2 (.I(_4535_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4957__A1 (.I(_4531_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4957__C (.I(_4231_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4958__I (.I(_4221_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4959__A2 (.I(_4527_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4959__B (.I(_4537_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4960__A2 (.I(_4514_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4961__I (.I(_4383_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4962__I (.I(_4541_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4964__A1 (.I(_4422_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4964__A2 (.I(_4194_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4965__A1 (.I(_4206_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4965__A2 (.I(_4543_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4965__A3 (.I(_4544_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4966__I (.I(_4545_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4967__I (.I(_4546_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4968__A1 (.I(_4542_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4968__A2 (.I(_4547_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4969__A3 (.I(_4548_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4970__I (.I(_4232_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4971__I (.I(_4550_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4972__A1 (.I(_4551_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4972__A2 (.I(_4242_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4972__A3 (.I(_4246_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4973__A1 (.I(_4154_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4975__A2 (.I(_4513_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4975__C (.I(_0285_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4977__A1 (.I(_4305_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4977__A2 (.I(_4306_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4977__A3 (.I(_0287_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4978__A1 (.I(_4348_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4978__A3 (.I(_4506_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4978__A4 (.I(_4509_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4979__I (.I(_4508_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4980__A1 (.I(_4348_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4980__B1 (.I(_4506_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4980__B2 (.I(_0290_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4981__A1 (.I(_0289_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4981__A2 (.I(_0291_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4982__A2 (.I(_0292_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4983__I (.I(_4248_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4984__A1 (.I(_0294_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4984__A2 (.I(_4261_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4985__I (.I(_0295_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4986__I (.I(\as2650.holding_reg[1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4987__A1 (.I(_4257_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4987__A2 (.I(_4386_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4988__A1 (.I(_0297_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4988__A2 (.I(_4332_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4989__A1 (.I(_4279_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4990__A1 (.I(_4381_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4990__A2 (.I(_4385_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4991__A1 (.I(\as2650.holding_reg[1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4991__A2 (.I(_0301_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4993__A1 (.I(\as2650.holding_reg[1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4993__A2 (.I(_0301_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4995__A3 (.I(_4302_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4996__B (.I(_4310_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4997__A2 (.I(_0307_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4998__A1 (.I(_4315_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4999__A1 (.I(_4302_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5000__A1 (.I(_4302_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5001__A1 (.I(_0310_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5001__B (.I(_4325_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5002__A1 (.I(_4277_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5002__A2 (.I(_4329_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5004__A1 (.I(_0297_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5005__A1 (.I(_4332_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5005__A2 (.I(_4386_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5005__B (.I(_4324_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5006__A3 (.I(_0313_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5007__A1 (.I(_4330_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5007__B (.I(_4338_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5008__A1 (.I(_4338_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5009__A2 (.I(_0319_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5011__A1 (.I(_0296_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5011__A2 (.I(_0321_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5014__A2 (.I(_4481_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5014__B1 (.I(_4460_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5014__C1 (.I(_0324_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5015__I (.I(_4478_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5016__A1 (.I(_4453_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5017__I (.I(_0327_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5018__I (.I(_0328_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5019__A1 (.I(\as2650.stack[7][9] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5020__A2 (.I(_4452_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5020__B (.I(_4454_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5021__A2 (.I(_4460_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5022__A1 (.I(\as2650.stack[0][9] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5022__A2 (.I(_4465_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5022__B1 (.I(_0324_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5025__A2 (.I(_0335_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5026__I (.I(_4542_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5027__A1 (.I(_4420_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5027__A2 (.I(_4488_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5028__I (.I(_0338_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5029__A1 (.I(_4277_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5029__A2 (.I(_4423_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5030__A1 (.I(_0339_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5030__A2 (.I(_0340_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5031__I (.I(_0341_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5032__I (.I(_0342_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5033__A1 (.I(_0337_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5034__A1 (.I(_4494_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5035__A2 (.I(_0323_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5035__B (.I(_0345_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5037__I (.I(\as2650.r123[0][2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5038__I (.I(_0287_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5039__A1 (.I(_4518_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5039__A2 (.I(_4523_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5040__A2 (.I(_4509_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5041__A1 (.I(_0348_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5041__A2 (.I(_0350_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5043__A1 (.I(_0352_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5043__A2 (.I(_0287_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5046__A2 (.I(_4505_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5047__A2 (.I(_0355_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5047__B1 (.I(_0356_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5047__B2 (.I(_0352_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5049__I (.I(_4520_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5050__I (.I(_0359_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5051__I (.I(_0360_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5052__I (.I(\as2650.r0[3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5053__I (.I(_0362_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5054__I (.I(_0363_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5055__A1 (.I(_0364_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5056__S (.I(_4516_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5057__I1 (.I(\as2650.r123[0][3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5057__I3 (.I(\as2650.r123_2[0][3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5057__S0 (.I(_4139_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5057__S1 (.I(_4516_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5058__A2 (.I(_0366_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5058__B1 (.I(_0367_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5058__B2 (.I(_4521_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5059__A1 (.I(_0365_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5059__A2 (.I(_0368_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5061__I (.I(_0370_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5062__I (.I(_0371_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5063__I (.I(net8));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5064__I (.I(_0373_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5065__I (.I(_0374_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5066__I (.I(_0375_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5067__A1 (.I(_4218_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5067__A2 (.I(_4507_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5067__B1 (.I(_4510_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5067__B2 (.I(_4533_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5068__A1 (.I(_4525_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5069__A1 (.I(_4399_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5069__A2 (.I(_0378_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5070__A1 (.I(_0376_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5071__A1 (.I(_4378_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5071__A2 (.I(_0372_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5072__A2 (.I(_4388_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5073__A1 (.I(_0361_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5073__B (.I(_4408_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5074__I (.I(_4503_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5075__A1 (.I(_0384_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5075__A2 (.I(_0350_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5076__A1 (.I(_4357_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5077__A1 (.I(_4359_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5077__A2 (.I(_4525_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5078__A1 (.I(_0386_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5078__A2 (.I(_0356_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5080__A1 (.I(_4354_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5080__A2 (.I(_0389_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5081__B (.I(_4345_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5082__A2 (.I(_0358_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5083__I (.I(_4312_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5084__I (.I(_4278_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5085__A1 (.I(_0393_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5085__A2 (.I(_0394_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5086__I (.I(_0395_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5087__I (.I(_4341_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5088__A1 (.I(\as2650.holding_reg[2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5088__A2 (.I(_0355_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5089__A1 (.I(\as2650.holding_reg[2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5089__A2 (.I(_0355_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5091__A1 (.I(\as2650.holding_reg[2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5091__A2 (.I(_0400_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5094__A1 (.I(_0297_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5095__A1 (.I(_0403_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5095__A2 (.I(_0307_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5096__A2 (.I(_0405_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5099__A2 (.I(_0310_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5099__B (.I(_0408_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5100__A2 (.I(_0310_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5100__A3 (.I(_0408_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5101__A1 (.I(_4277_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5101__A2 (.I(_4324_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5102__B (.I(_0411_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5103__I (.I(\as2650.holding_reg[2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5105__A2 (.I(_4526_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5106__A1 (.I(_0413_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5106__B (.I(_4314_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5107__A1 (.I(_4315_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5108__I (.I(_4330_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5109__A1 (.I(_0397_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5109__A2 (.I(_0398_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5109__B2 (.I(_0313_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5109__C2 (.I(_0418_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5110__A1 (.I(_0395_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5110__A2 (.I(_0408_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5111__A1 (.I(_0396_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5111__A2 (.I(_0419_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5112__I (.I(_0421_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5113__A2 (.I(_0422_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5115__A2 (.I(_4452_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5115__B (.I(_4454_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5117__I (.I(_0426_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5118__A1 (.I(\as2650.stack[2][10] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5118__A2 (.I(_0427_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5119__I (.I(_4465_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5120__I (.I(_4469_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5121__A1 (.I(\as2650.stack[0][10] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5121__A2 (.I(_0429_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5121__B1 (.I(_0430_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5123__A2 (.I(_0429_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5123__B1 (.I(_4470_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5124__B1 (.I(_0427_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5124__B2 (.I(\as2650.stack[6][10] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5125__A1 (.I(_4477_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5126__A2 (.I(_0435_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5127__A1 (.I(_0361_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5127__A2 (.I(_0342_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5129__A2 (.I(_0436_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5130__A2 (.I(_0424_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5132__I (.I(\as2650.r123[0][3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5133__A1 (.I(\as2650.holding_reg[3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5133__A2 (.I(_0370_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5134__A1 (.I(\as2650.holding_reg[3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5134__A2 (.I(_0371_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5135__A1 (.I(_0442_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5137__A1 (.I(_0395_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5138__I (.I(_0393_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5139__A1 (.I(_0447_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5139__A2 (.I(_4314_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5141__A1 (.I(_4257_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5141__A2 (.I(_4525_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5142__A1 (.I(_0413_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5143__A1 (.I(_0398_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5143__A2 (.I(_0451_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5144__A2 (.I(_0405_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5146__A1 (.I(_0448_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5146__A2 (.I(_0454_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5147__A2 (.I(_4522_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5148__A1 (.I(_0359_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5148__A2 (.I(_4142_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5149__A1 (.I(_4518_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5149__A2 (.I(_0457_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5150__A1 (.I(_0413_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5150__A2 (.I(_0456_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5150__B2 (.I(_0310_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5150__B3 (.I(_0398_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5152__I (.I(\as2650.holding_reg[3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5153__A1 (.I(_0365_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5153__A2 (.I(_0368_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5156__A2 (.I(_0464_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5157__A1 (.I(_0461_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5159__A1 (.I(_0393_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5159__A2 (.I(_0467_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5160__I (.I(_4191_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5161__A1 (.I(_0469_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5161__A2 (.I(_0464_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5162__A1 (.I(_0461_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5162__A2 (.I(_4422_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5162__B (.I(_4336_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5163__A1 (.I(_0411_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5163__A2 (.I(_0460_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5163__B2 (.I(_4225_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5164__I (.I(_4279_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5165__A1 (.I(_0397_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5165__A2 (.I(_0442_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5165__C (.I(_0473_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5166__A1 (.I(_0446_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5166__A2 (.I(_0474_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5168__A2 (.I(_4505_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5169__A1 (.I(_4304_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5169__A2 (.I(_4386_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5169__A3 (.I(_4524_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5170__A1 (.I(_0477_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5170__A2 (.I(_0478_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5170__B (.I(_0352_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5171__A1 (.I(_4518_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5171__A2 (.I(_4523_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5171__A3 (.I(_0365_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5171__A4 (.I(_0368_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5173__A1 (.I(_4509_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5173__A2 (.I(_0481_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5174__A1 (.I(_4524_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5174__A2 (.I(_0290_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5175__A1 (.I(_0348_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5175__B2 (.I(_0370_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5177__I (.I(_4269_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5178__I (.I(_4359_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5179__A1 (.I(_0477_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5179__A2 (.I(_0478_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5180__A1 (.I(_0384_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5181__A1 (.I(_0487_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5181__A2 (.I(_0464_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5182__I (.I(_0490_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5183__I (.I(_0364_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5184__I (.I(_4379_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5185__I1 (.I(\as2650.r123[0][4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5185__I3 (.I(\as2650.r123_2[0][4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5185__S0 (.I(_4196_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5185__S1 (.I(_0493_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5186__A1 (.I(_4521_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5186__A2 (.I(_0494_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5187__S (.I(_4516_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5188__A2 (.I(_0496_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5189__I (.I(\as2650.r0[4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5190__I (.I(_0498_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5191__I (.I(_0499_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5192__A1 (.I(_0500_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5193__A1 (.I(_0495_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5193__A3 (.I(_0501_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5194__I (.I(_0502_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5195__I (.I(_0503_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5196__I (.I(_0504_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5197__I (.I(net9));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5198__I (.I(_0506_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5199__I (.I(_0507_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5200__A1 (.I(_4218_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5200__A2 (.I(_0355_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5200__A3 (.I(_4507_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5201__A1 (.I(_4533_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5201__A2 (.I(_4524_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5201__A3 (.I(_4510_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5204__A1 (.I(_4396_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5204__A2 (.I(_0512_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5205__A1 (.I(_0508_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5205__A2 (.I(_4399_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5206__A2 (.I(_0505_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5206__C (.I(_4221_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5207__I (.I(_4220_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5208__A1 (.I(_4212_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5208__A2 (.I(_0516_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5209__A1 (.I(_0517_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5209__A2 (.I(_4526_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5209__B (.I(_4545_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5210__A1 (.I(_0492_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5210__A2 (.I(_4545_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5211__A1 (.I(_4269_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5212__A1 (.I(_0486_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5212__A2 (.I(_0491_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5212__C (.I(_4247_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5213__A1 (.I(_4345_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5213__A2 (.I(_0485_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5213__C (.I(_4262_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5214__A2 (.I(_0476_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5215__I (.I(_0523_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5216__I (.I(_0328_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5217__I (.I(_0525_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5218__I (.I(_0426_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5219__A2 (.I(_4450_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5219__B1 (.I(_4469_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5221__A1 (.I(\as2650.stack[0][11] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5221__A2 (.I(_0429_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5221__B1 (.I(_0527_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5221__B2 (.I(\as2650.stack[2][11] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5222__A2 (.I(_0429_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5222__B1 (.I(_0430_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5223__A2 (.I(_4478_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5223__B1 (.I(_0527_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5223__B2 (.I(\as2650.stack[6][11] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5224__A1 (.I(_0526_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5225__A2 (.I(_0533_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5226__I (.I(_0492_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5227__A1 (.I(_0535_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5228__A1 (.I(_4494_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5230__A2 (.I(_0524_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5230__B (.I(_0537_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5232__I (.I(\as2650.r123[0][4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5233__A1 (.I(_0495_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5233__A3 (.I(_0501_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5234__I (.I(_0541_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5235__A2 (.I(_0542_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5236__I (.I(_4325_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5237__A1 (.I(_0461_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5237__A2 (.I(_0371_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5239__A1 (.I(_0543_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5242__I (.I(_4332_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5243__A1 (.I(_0549_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5243__A2 (.I(_0550_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5244__A1 (.I(_0548_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5244__A2 (.I(_0504_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5245__I (.I(_4336_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5246__A1 (.I(_0544_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5246__B2 (.I(_0553_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5247__I (.I(_4315_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5248__A1 (.I(_0549_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5248__A2 (.I(_0504_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5249__B2 (.I(_0442_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5251__A1 (.I(_0549_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5252__A1 (.I(_4488_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5252__A2 (.I(_0504_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5253__I (.I(_0560_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5254__I (.I(_4338_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5255__A1 (.I(_0555_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5255__B1 (.I(_0561_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5255__B2 (.I(_0418_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5255__C (.I(_0562_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5257__I (.I(_0562_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5258__I (.I(_0542_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5259__A2 (.I(_0566_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5260__A1 (.I(_0565_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5260__B (.I(_0396_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5261__A1 (.I(_0396_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5261__A2 (.I(_0543_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5262__I (.I(_0569_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5264__A1 (.I(_0477_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5264__A2 (.I(_0541_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5265__A1 (.I(_4359_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5265__A2 (.I(_0503_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5266__A1 (.I(_0290_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5266__A2 (.I(_0481_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5266__A3 (.I(_0502_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5267__A1 (.I(_0290_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5267__A2 (.I(_0481_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5267__B (.I(_0502_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5268__A1 (.I(_0384_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5269__A1 (.I(_0571_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5270__I (.I(_0577_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5271__I (.I(_0500_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5272__I (.I(_0579_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5273__I1 (.I(\as2650.r123[0][5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5273__I3 (.I(\as2650.r123_2[0][5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5273__S0 (.I(_4196_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5273__S1 (.I(_0493_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5274__A1 (.I(_4521_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5274__A2 (.I(_0581_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5275__S (.I(_0493_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5276__A2 (.I(_0583_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5277__I (.I(\as2650.r0[5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5278__I (.I(_0585_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5279__A1 (.I(_0586_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5280__A3 (.I(_0587_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5281__I (.I(_0588_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5284__I (.I(_0591_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5285__I (.I(_0592_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5286__I (.I(net10));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5287__I (.I(_0594_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5288__I (.I(_0595_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5289__I (.I(_0596_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5290__I (.I(_4396_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5291__A1 (.I(_4508_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5293__A1 (.I(_4155_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5293__A2 (.I(_0600_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5294__B1 (.I(_0599_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5294__B2 (.I(_0601_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5295__A1 (.I(_0503_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5296__A2 (.I(_0603_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5297__A1 (.I(_0597_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5297__A2 (.I(_0598_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5298__A1 (.I(_4378_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5298__A2 (.I(_0593_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5299__A2 (.I(_0372_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5300__A1 (.I(_0580_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5301__A2 (.I(_0578_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5301__C (.I(_0285_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5303__I (.I(_4348_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5304__A1 (.I(_0348_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5305__A1 (.I(_0610_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5305__A2 (.I(_0503_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5305__B2 (.I(_0611_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5306__I (.I(_0613_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5307__A2 (.I(_0614_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5308__A2 (.I(_0570_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5309__I (.I(_0580_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5310__I (.I(_4426_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5313__I (.I(_0620_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5314__I (.I(_4452_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5315__A2 (.I(_0622_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5315__B (.I(_4454_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5316__I (.I(_4460_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5317__A1 (.I(\as2650.stack[2][12] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5317__A2 (.I(_0624_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5318__I (.I(_0324_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5319__A1 (.I(\as2650.stack[0][12] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5319__A2 (.I(_4482_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5319__B1 (.I(_0626_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5319__B2 (.I(\as2650.stack[1][12] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5321__A2 (.I(_4482_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5321__B1 (.I(_0626_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5322__A2 (.I(_4479_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5322__B1 (.I(_4461_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5323__A1 (.I(_4477_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5324__A2 (.I(_0631_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5325__A1 (.I(_0617_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5325__A2 (.I(_0621_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5325__B2 (.I(_0632_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5326__A2 (.I(_0616_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5326__B (.I(_0633_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5327__A1 (.I(_0540_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5328__I (.I(\as2650.r123[0][5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5329__I (.I(_0395_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5331__A3 (.I(_0587_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5332__I (.I(_0638_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5333__A1 (.I(_0637_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5333__A2 (.I(_0639_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5335__A2 (.I(_0591_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5337__A1 (.I(_0543_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5339__A1 (.I(_0544_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5340__B1 (.I(_0560_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5341__A1 (.I(_0641_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5341__A2 (.I(_0647_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5342__A2 (.I(_0647_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5343__A1 (.I(_0555_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5344__I (.I(_0418_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5345__A2 (.I(_4191_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5346__A2 (.I(_0591_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5348__A1 (.I(_0637_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5348__A2 (.I(_0548_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5349__A1 (.I(_0654_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5349__A2 (.I(_0592_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5350__A1 (.I(_0651_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5350__A2 (.I(_0653_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5350__B2 (.I(_0553_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5350__C (.I(_0562_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5352__A1 (.I(_0637_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5352__A2 (.I(_0638_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5353__A1 (.I(_0565_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5353__B (.I(_0396_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5354__A1 (.I(_0636_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5354__A2 (.I(_0641_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5355__I (.I(_0661_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5357__A2 (.I(_4505_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5357__A4 (.I(_0541_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5358__A2 (.I(_0664_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5359__A1 (.I(_0611_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5360__A1 (.I(_0610_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5360__B2 (.I(_4350_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5361__I (.I(_0667_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5362__I (.I(_0586_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5363__I (.I(_0669_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5364__I (.I(\as2650.r0[6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5365__I (.I(_0671_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5366__A1 (.I(_0672_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5366__A2 (.I(_4142_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5367__S (.I(_0493_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5368__A1 (.I(_4369_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5368__A2 (.I(_0674_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5369__I1 (.I(\as2650.r123[0][6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5369__I3 (.I(\as2650.r123_2[0][6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5369__S0 (.I(_4196_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5369__S1 (.I(_4148_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5370__A2 (.I(_0676_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5371__A1 (.I(_0673_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5372__I (.I(_0678_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5373__I (.I(_0679_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5374__I (.I(_0680_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5375__I (.I(net1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5376__I (.I(_0682_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5377__I (.I(_0683_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5378__I (.I(_0684_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5379__A2 (.I(_4506_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5379__A3 (.I(_0370_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5379__A4 (.I(_0542_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5380__A2 (.I(_4193_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5381__A1 (.I(_4155_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5381__A2 (.I(_0687_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5382__A1 (.I(_0601_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5382__A2 (.I(_0599_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5382__A3 (.I(_0542_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5382__B1 (.I(_0686_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5382__B2 (.I(_0688_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5384__A1 (.I(_0598_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5384__A2 (.I(_0690_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5385__A1 (.I(_0685_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5385__C (.I(_4378_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5386__A2 (.I(_0681_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5387__I (.I(_0505_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5388__A1 (.I(_0517_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5388__A2 (.I(_0694_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5388__B (.I(_4546_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5389__A1 (.I(_0670_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5389__A2 (.I(_4547_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5389__B1 (.I(_0693_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5390__A1 (.I(_0571_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5390__C1 (.I(_0487_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5390__C2 (.I(_0591_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5391__I (.I(_0697_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5392__A1 (.I(_0486_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5392__A2 (.I(_0698_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5394__A1 (.I(_4354_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5394__C (.I(_0700_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5395__A1 (.I(_0285_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5395__A2 (.I(_0668_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5395__C (.I(_0295_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5396__A1 (.I(_0296_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5396__A2 (.I(_0662_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5397__A1 (.I(\as2650.stack[7][13] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5397__B1 (.I(_4466_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5397__B2 (.I(\as2650.stack[4][13] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5397__C1 (.I(\as2650.stack[5][13] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5397__C2 (.I(_4470_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5398__A1 (.I(\as2650.stack[6][13] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5398__A2 (.I(_4461_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5399__A2 (.I(_4481_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5399__B1 (.I(_0324_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5401__A1 (.I(\as2650.stack[3][13] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5401__A2 (.I(_4479_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5401__B1 (.I(_0427_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5401__B2 (.I(\as2650.stack[2][13] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5401__C (.I(_0707_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5402__B2 (.I(_0526_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5403__A2 (.I(_0709_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5404__I (.I(_0670_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5405__A1 (.I(_0711_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5407__A1 (.I(_4274_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5407__A2 (.I(_0703_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5407__B (.I(_0713_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5409__I (.I(\as2650.r123[0][6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5410__A1 (.I(_0673_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5411__I (.I(_0716_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5413__A2 (.I(_0718_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5414__I (.I(_0719_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5415__I (.I(_0719_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5416__A2 (.I(_0653_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5417__A2 (.I(_0647_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5419__A2 (.I(_0720_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5420__A1 (.I(_0555_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5420__A2 (.I(_0724_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5422__A1 (.I(_0719_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5422__A2 (.I(_0727_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5422__B (.I(_0411_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5423__A1 (.I(_0720_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5423__A2 (.I(_0727_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5425__A2 (.I(_0469_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5426__A1 (.I(_4427_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5426__A2 (.I(_0679_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5427__A2 (.I(_0548_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5428__A1 (.I(_0654_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5428__A2 (.I(_0680_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5429__A1 (.I(_0651_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5429__A2 (.I(_0732_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5429__B2 (.I(_0553_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5429__C (.I(_0562_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5431__A2 (.I(_0718_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5432__A1 (.I(_0565_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5432__A2 (.I(_0737_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5432__B (.I(_0636_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5433__A1 (.I(_0636_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5433__A2 (.I(_0720_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5435__A1 (.I(_0638_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5435__A2 (.I(_0664_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5435__A3 (.I(_0716_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5436__A2 (.I(_0686_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5436__B (.I(_0678_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5438__A1 (.I(_0502_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5438__A2 (.I(_0588_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5439__A1 (.I(_0599_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5440__A1 (.I(_0745_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5440__A2 (.I(_0716_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5441__A1 (.I(_0348_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5442__A1 (.I(_0610_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5442__A2 (.I(_0678_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5442__B2 (.I(_0611_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5443__I (.I(_0748_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5444__I (.I(_0672_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5445__I (.I(_0750_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5446__I (.I(_0751_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5447__I (.I(_4376_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5448__I (.I(_0753_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5449__I (.I(net2));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5451__I (.I(_0756_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5452__I (.I(_0757_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5453__I (.I(_0758_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5454__A1 (.I(_4533_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5455__A1 (.I(_4218_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5455__A2 (.I(_0638_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5455__A3 (.I(_0664_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5456__A1 (.I(_0760_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5457__A1 (.I(_0679_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5458__A1 (.I(_0598_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5458__A2 (.I(_0763_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5459__A1 (.I(_0759_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5459__C (.I(_4231_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5460__A2 (.I(_0754_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5461__A1 (.I(_0517_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5461__A2 (.I(_0593_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5461__B (.I(_4546_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5462__A1 (.I(_0752_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5462__A2 (.I(_4547_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5462__B1 (.I(_0766_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5463__A1 (.I(_0384_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5464__A1 (.I(_0487_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5464__A2 (.I(_0679_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5464__B2 (.I(_0571_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5465__I (.I(_0770_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5466__A1 (.I(_0486_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5466__A2 (.I(_0771_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5467__A1 (.I(_4354_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5467__C (.I(_0700_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5468__A1 (.I(_0285_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5468__A2 (.I(_0749_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5468__C (.I(_0295_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5469__A1 (.I(_0296_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5469__A2 (.I(_0740_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5470__B1 (.I(_0527_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5470__B2 (.I(\as2650.stack[6][14] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5471__A1 (.I(\as2650.stack[4][14] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5471__A2 (.I(_4481_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5471__B1 (.I(_0430_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5471__B2 (.I(\as2650.stack[5][14] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5472__A2 (.I(_4465_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5472__B1 (.I(_4469_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5474__A1 (.I(\as2650.stack[3][14] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5474__A2 (.I(_4478_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5474__B1 (.I(_0527_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5474__C (.I(_0779_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5475__B2 (.I(_0526_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5476__A1 (.I(_4445_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5476__A2 (.I(_0781_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5477__A1 (.I(_0752_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5479__A1 (.I(_4274_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5479__A2 (.I(_0775_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5479__B (.I(_0784_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5481__I (.I(\as2650.r123[0][7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5482__I (.I(_4494_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5483__I (.I(_4367_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5484__I (.I(_0788_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5485__I (.I(_0789_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5486__I (.I(_0790_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5487__A1 (.I(_0791_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5487__A2 (.I(_0620_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5489__A2 (.I(_4376_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5490__I (.I(_0794_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5492__A1 (.I(_0737_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5492__A2 (.I(_0732_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5494__A1 (.I(_4368_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5495__A2 (.I(_0799_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5497__B (.I(_0801_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5498__A1 (.I(_0724_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5498__A2 (.I(_0794_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5499__B (.I(_0448_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5500__I (.I(_0737_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5501__A1 (.I(_0719_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5501__A2 (.I(_0727_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5502__A1 (.I(_0794_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5503__A1 (.I(_0544_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5504__A2 (.I(_0550_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5505__A1 (.I(_0550_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5505__A2 (.I(_4376_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5506__A1 (.I(_4336_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5507__A1 (.I(_0313_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5509__I (.I(_0447_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5510__A2 (.I(_0799_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5510__B (.I(_0814_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5511__A1 (.I(_0651_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5511__A2 (.I(_0815_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5513__I (.I(_0799_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5514__A2 (.I(_0565_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5514__A3 (.I(_0818_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5515__A1 (.I(_0473_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5516__A1 (.I(_0636_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5516__A2 (.I(_0795_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5517__A1 (.I(_0799_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5518__A1 (.I(_0611_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5519__A1 (.I(_0599_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5520__A1 (.I(_4374_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5520__A2 (.I(_0824_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5521__A1 (.I(_4375_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5521__A2 (.I(_0610_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5521__B1 (.I(_0825_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5521__B2 (.I(_4350_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5523__I (.I(_0827_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5524__A1 (.I(_4375_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5524__A2 (.I(_0487_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5524__B2 (.I(_0571_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5524__C1 (.I(_0825_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5525__I (.I(_0829_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5526__A1 (.I(_4408_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5526__A2 (.I(_0830_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5526__B (.I(_0700_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5527__I0 (.I(_0760_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5528__A1 (.I(_4375_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5529__I (.I(_0833_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5530__I (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5532__I (.I(_0836_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5533__A1 (.I(_0837_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5533__A2 (.I(_0598_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5533__B (.I(_4231_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5534__A2 (.I(_0834_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5535__A1 (.I(_4320_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5535__A2 (.I(_4334_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5535__B (.I(_4321_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5536__A2 (.I(_0840_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5538__A1 (.I(_0517_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5538__A2 (.I(_0681_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5538__B (.I(_4546_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5539__A1 (.I(_0790_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5539__A2 (.I(_4547_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5539__B1 (.I(_0842_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5539__C (.I(_0486_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5540__A1 (.I(_0700_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5540__A2 (.I(_0828_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5540__C (.I(_0295_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5541__A1 (.I(_0296_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5541__A2 (.I(_0821_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5542__A2 (.I(_0846_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5544__I (.I(_4295_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5546__I (.I(_0849_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5547__I (.I(_0850_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5548__I (.I(_4204_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5550__A1 (.I(_4488_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5551__A1 (.I(_0853_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5551__A2 (.I(_0854_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5552__A1 (.I(_0852_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5552__A2 (.I(_0855_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5553__I (.I(_0856_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5555__A2 (.I(_0626_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5555__A3 (.I(_0858_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5556__I (.I(_0859_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5557__I (.I(_0860_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5558__I (.I(\as2650.pc[0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5559__I (.I(_0862_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5560__I (.I(_0863_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5561__I (.I(_0864_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5562__I (.I(_0850_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5563__I (.I(_4214_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5564__I (.I(_4215_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5565__A2 (.I(_4369_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5565__A3 (.I(_4313_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5566__A1 (.I(_4255_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5566__A2 (.I(_0869_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5567__I (.I(_0870_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5568__A1 (.I(_0868_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5568__A2 (.I(_0871_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5569__A1 (.I(_0867_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5569__A2 (.I(_0872_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5570__I (.I(_4184_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5571__A2 (.I(_4193_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5572__I (.I(_4180_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5573__I (.I(_0876_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5574__A2 (.I(_4175_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5575__I (.I(_0878_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5576__A1 (.I(_0877_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5576__A2 (.I(_0879_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5577__I (.I(\as2650.addr_buff[7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5578__I (.I(_4254_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5579__I (.I(_4208_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5580__I (.I(\as2650.cycle[1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5581__I (.I(_4238_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5583__A2 (.I(_0885_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5584__A3 (.I(_0884_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5585__A1 (.I(_0883_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5586__A1 (.I(_0881_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5586__A2 (.I(_0882_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5586__B (.I(_0889_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5587__A1 (.I(_0877_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5587__A2 (.I(_0870_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5588__A1 (.I(_0836_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5588__B1 (.I(_0890_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5588__B2 (.I(_0891_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5590__A1 (.I(_0893_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5590__A3 (.I(_4172_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5591__A1 (.I(_0884_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5591__A2 (.I(_4208_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5592__I (.I(_0895_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5593__A1 (.I(_0447_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5593__A2 (.I(_0896_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5594__I (.I(_0891_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5595__A1 (.I(_0873_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5595__A2 (.I(_0875_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5595__A3 (.I(_0892_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5595__B1 (.I(_0897_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5595__B2 (.I(_0898_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5596__A1 (.I(_4152_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5596__A2 (.I(_0899_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5597__I (.I(_0900_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5598__A1 (.I(_0866_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5598__A2 (.I(_4466_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5598__A3 (.I(_0901_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5599__I (.I(_0902_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5600__I (.I(_0902_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5601__A1 (.I(\as2650.stack[5][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5602__A1 (.I(_0865_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5602__A2 (.I(_0903_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5604__A1 (.I(_0848_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5605__I (.I(_0337_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5607__I (.I(_0909_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5608__I (.I(_0910_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5609__I (.I(_0911_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5610__I (.I(_0902_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5611__I0 (.I(_0912_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5611__I1 (.I(\as2650.stack[5][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5611__S (.I(_0913_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5612__I (.I(_0859_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5613__I0 (.I(_0908_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5613__S (.I(_0915_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5615__I (.I(_0361_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5616__I (.I(_0917_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5617__I (.I(\as2650.pc[2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5618__I (.I(_0919_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5620__I0 (.I(_0921_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5620__I1 (.I(\as2650.stack[5][2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5620__S (.I(_0913_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5621__I0 (.I(_0918_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5621__S (.I(_0915_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5623__I (.I(_0535_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5624__I (.I(_0924_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5626__I (.I(_0926_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5628__A1 (.I(\as2650.stack[5][3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5629__A1 (.I(_0928_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5629__A2 (.I(_0903_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5630__I0 (.I(_0925_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5630__S (.I(_0860_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5632__I (.I(_0617_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5634__A1 (.I(\as2650.stack[5][4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5634__A2 (.I(_0913_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5635__A1 (.I(_0933_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5635__A2 (.I(_0903_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5636__A1 (.I(_0915_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5637__A1 (.I(_0932_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5638__I (.I(_0711_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5641__I (.I(_0939_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5642__A1 (.I(\as2650.stack[5][5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5642__A2 (.I(_0913_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5643__A1 (.I(_0940_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5644__A1 (.I(_0915_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5645__A1 (.I(_0938_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5646__I (.I(_0752_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5647__I (.I(\as2650.pc[6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5648__I (.I(_0945_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5649__I (.I(_0946_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5650__I (.I(_0947_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5651__I0 (.I(_0948_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5651__I1 (.I(\as2650.stack[5][6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5651__S (.I(_0902_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5652__I0 (.I(_0944_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5652__S (.I(_0860_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5654__I (.I(_0791_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5655__I (.I(\as2650.pc[7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5657__A1 (.I(\as2650.stack[5][7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5658__A1 (.I(_0953_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5658__A2 (.I(_0903_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5659__I0 (.I(_0951_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5659__S (.I(_0860_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5661__I (.I(_0850_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5662__A1 (.I(_0957_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5662__A2 (.I(_0430_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5663__A1 (.I(_0856_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5663__A2 (.I(_0900_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5665__A2 (.I(_0960_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5666__I (.I(_0961_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5667__I (.I(_0962_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5668__I (.I(\as2650.pc[8] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5672__I (.I(_0967_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5673__I (.I(_4152_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5674__A2 (.I(_0854_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5675__I (.I(_0970_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5676__A1 (.I(_0294_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5676__A3 (.I(_0971_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5677__I (.I(_0972_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5678__A1 (.I(\as2650.r123[0][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5678__A2 (.I(_4153_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5678__A3 (.I(_0855_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5679__A1 (.I(_0966_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5679__A2 (.I(_0968_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5679__B2 (.I(\as2650.r123_2[0][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5679__C (.I(_0974_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5680__I (.I(_0975_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5681__I (.I(_0962_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5683__A1 (.I(_0963_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5683__A2 (.I(_0976_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5685__I (.I(_0967_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5686__I (.I(_4415_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5687__I (.I(_0971_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5688__A2 (.I(_0981_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5689__A1 (.I(_0979_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5689__B2 (.I(\as2650.r123_2[0][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5689__C (.I(_0983_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5690__I (.I(_0984_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5691__I (.I(_0961_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5692__A2 (.I(_0986_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5693__A1 (.I(_0963_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5693__A2 (.I(_0985_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5696__I (.I(_0989_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5697__A2 (.I(_0981_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5698__A1 (.I(_0990_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5698__B2 (.I(\as2650.r123_2[0][2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5698__C (.I(_0991_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5699__I (.I(_0992_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5700__A1 (.I(\as2650.stack[6][10] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5700__A2 (.I(_0986_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5701__A1 (.I(_0963_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5701__A2 (.I(_0993_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5702__I (.I(\as2650.pc[11] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5703__I (.I(_0995_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5705__A2 (.I(_0981_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5706__A1 (.I(_0997_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5706__B2 (.I(\as2650.r123_2[0][3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5706__C (.I(_0998_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5707__I (.I(_0999_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5708__A1 (.I(\as2650.stack[6][11] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5708__A2 (.I(_0986_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5709__A1 (.I(_0963_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5709__A2 (.I(_1000_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5710__I (.I(\as2650.pc[12] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5712__A1 (.I(_0540_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5713__A1 (.I(_1003_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5713__B1 (.I(_0972_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5713__B2 (.I(\as2650.r123_2[0][4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5713__C (.I(_1004_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5714__I (.I(_1005_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5715__A2 (.I(_0986_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5716__A2 (.I(_1006_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5718__I (.I(_0971_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5719__A3 (.I(_1009_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5720__A1 (.I(_1008_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5720__A2 (.I(_0858_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5720__B1 (.I(_0972_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5720__B2 (.I(\as2650.r123_2[0][5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5720__C (.I(_1010_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5721__I (.I(_1011_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5722__A1 (.I(\as2650.stack[6][13] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5722__A2 (.I(_0962_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5723__A2 (.I(_1012_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5724__A3 (.I(_1009_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5725__A1 (.I(\as2650.pc[14] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5725__A2 (.I(_0858_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5725__B1 (.I(_0972_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5725__B2 (.I(\as2650.r123_2[0][6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5725__C (.I(_1014_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5727__A1 (.I(\as2650.stack[6][14] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5727__A2 (.I(_0962_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5728__A2 (.I(_1016_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5729__A1 (.I(_0866_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5729__A2 (.I(_4466_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5731__A2 (.I(_1019_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5733__I (.I(_1021_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5734__I (.I(_1021_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5736__A1 (.I(_0976_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5736__A2 (.I(_1022_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5738__A2 (.I(_1025_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5739__A1 (.I(_0985_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5739__A2 (.I(_1022_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5740__A2 (.I(_1025_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5741__A1 (.I(_0993_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5741__A2 (.I(_1022_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5742__A2 (.I(_1025_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5743__A1 (.I(_1000_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5743__A2 (.I(_1022_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5744__A2 (.I(_1025_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5745__A1 (.I(_1006_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5746__A1 (.I(\as2650.stack[5][13] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5746__A2 (.I(_1021_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5747__A1 (.I(_1012_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5748__A1 (.I(\as2650.stack[5][14] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5748__A2 (.I(_1021_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5749__A1 (.I(_1016_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5750__I (.I(\as2650.r123_2[0][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5752__I (.I(_4200_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5753__A1 (.I(_1033_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5753__A2 (.I(_1034_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5754__A1 (.I(_4248_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5754__A2 (.I(_4151_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5755__A1 (.I(_4143_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5755__A2 (.I(_1036_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5756__A1 (.I(_4189_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5756__A2 (.I(_1037_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5757__A2 (.I(_1037_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5758__A2 (.I(_4198_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5758__A3 (.I(_4151_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5759__A1 (.I(_4157_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5759__A2 (.I(_4242_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5759__A3 (.I(_4245_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5759__A4 (.I(_1040_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5760__A1 (.I(_4210_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5760__A2 (.I(_1040_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5761__A1 (.I(_0876_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5761__A2 (.I(_0688_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5762__A1 (.I(_4180_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5762__A2 (.I(_4249_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5762__A3 (.I(_4341_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5763__A1 (.I(_1043_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5764__A1 (.I(_4223_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5764__A2 (.I(_1045_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5765__A2 (.I(_4261_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5766__A1 (.I(_4195_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5766__A2 (.I(_1042_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5767__A1 (.I(_1047_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5768__A1 (.I(_1042_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5768__A2 (.I(_1046_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5769__A2 (.I(_1039_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5769__A3 (.I(_1041_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5770__A2 (.I(_1051_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5771__A2 (.I(_1035_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5771__B (.I(_1052_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5771__C (.I(_4438_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5772__I (.I(_1053_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5774__I (.I(_1052_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5775__I (.I(_1041_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5776__I (.I(_1039_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5778__I (.I(_1041_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5779__I (.I(_1039_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5782__I (.I(_4377_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5783__A1 (.I(_4220_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5783__A2 (.I(_1042_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5785__A1 (.I(_4228_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5785__A2 (.I(_1042_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5786__I (.I(_1067_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5788__A1 (.I(_4395_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5788__A2 (.I(_1037_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5791__A1 (.I(_4398_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5792__A1 (.I(_4392_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5792__A2 (.I(_1071_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5792__C (.I(_1067_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5793__A1 (.I(_0301_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5795__A1 (.I(_1064_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5796__A1 (.I(_4406_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5797__A1 (.I(_1061_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5798__A1 (.I(_4361_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5798__A2 (.I(_1059_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5798__B (.I(_1060_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5799__A1 (.I(_4353_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5799__A2 (.I(_1057_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5799__B (.I(_1080_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5800__I (.I(_1047_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5801__I (.I(_1082_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5802__I0 (.I(_4344_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5803__A1 (.I(_4472_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5803__A2 (.I(_4484_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5804__I (.I(_4170_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5805__A1 (.I(_1086_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5805__A2 (.I(_0341_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5806__A1 (.I(_1087_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5806__A2 (.I(_1036_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5807__I (.I(_0294_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5808__A1 (.I(_1089_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5809__A1 (.I(_4295_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5809__A2 (.I(_0621_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5809__B1 (.I(_1085_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5810__A2 (.I(_1084_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5812__I (.I(\as2650.r123_2[0][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5813__A1 (.I(_1033_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5813__A2 (.I(_4261_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5814__I (.I(_4233_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5815__A1 (.I(_1095_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5815__A2 (.I(_4268_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5815__A3 (.I(_1040_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5816__I (.I(_1096_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5817__A1 (.I(_4513_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5819__I (.I(_4334_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5821__I (.I(_1067_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5823__I (.I(_4529_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5825__A1 (.I(_0301_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5825__A2 (.I(_4534_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5826__A1 (.I(_1106_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5826__A2 (.I(_1071_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5827__A1 (.I(_1104_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5828__A1 (.I(_0400_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5830__A1 (.I(_1100_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5830__C (.I(_1110_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5831__A1 (.I(_4542_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5831__C (.I(_1059_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5832__A1 (.I(_1060_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5832__A3 (.I(_1112_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5833__A1 (.I(_0292_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5833__A2 (.I(_1057_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5834__A1 (.I(_0321_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5834__A2 (.I(_1094_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5835__A1 (.I(_1094_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5838__A1 (.I(_1089_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5838__A2 (.I(_1118_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5838__A3 (.I(_4444_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5839__A1 (.I(_0335_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5839__A2 (.I(_1119_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5841__A2 (.I(_1116_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5843__I (.I(\as2650.r123_2[0][2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5844__I (.I(_1053_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5845__A1 (.I(_0436_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5846__I (.I(_1052_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5848__A1 (.I(_0378_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5848__A2 (.I(_1071_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5849__A1 (.I(_0376_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5850__A1 (.I(_0372_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5850__B (.I(_1127_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5851__A1 (.I(_4388_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5851__C (.I(_1110_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5852__A1 (.I(_0360_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5852__C (.I(_1061_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5853__A2 (.I(_1037_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5855__A1 (.I(_0389_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5855__B (.I(_1134_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5856__I (.I(_1041_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5857__A1 (.I(_0358_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5857__A2 (.I(_1136_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5858__A1 (.I(_1132_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5858__C (.I(_1094_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5859__A1 (.I(_0422_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5859__A2 (.I(_1094_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5860__A2 (.I(_1139_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5863__I (.I(\as2650.r123_2[0][3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5864__A1 (.I(_0533_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5864__A2 (.I(_1119_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5866__I (.I(_1082_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5867__A1 (.I(_4188_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5867__A2 (.I(_1040_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5868__I (.I(_0508_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5869__A1 (.I(_1147_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5869__A2 (.I(_1146_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5870__A1 (.I(_0512_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5870__A2 (.I(_1146_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5871__A1 (.I(_0566_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5871__B (.I(_1127_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5872__A1 (.I(_4527_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5872__C (.I(_1110_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5873__A1 (.I(_0535_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5873__C (.I(_1061_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5874__A1 (.I(_0491_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5874__B (.I(_1134_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5875__A1 (.I(_0485_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5875__A2 (.I(_1134_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5875__B1 (.I(_1152_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5876__A1 (.I(_0446_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5876__A2 (.I(_0474_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5876__B (.I(_1082_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5877__A1 (.I(_1145_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5877__B (.I(_1155_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5878__A2 (.I(_1156_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5881__I (.I(\as2650.r123_2[0][4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5883__A1 (.I(_0617_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5883__A2 (.I(_0621_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5883__B1 (.I(_0632_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5884__A1 (.I(_0603_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5885__I (.I(_4228_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5886__A1 (.I(_1033_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5886__A2 (.I(_4420_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5886__A3 (.I(_4204_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5886__A4 (.I(_4211_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5887__A1 (.I(_1163_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5887__A2 (.I(_1164_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5888__A1 (.I(_0596_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5888__C (.I(_1165_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5889__A1 (.I(_0592_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5890__A1 (.I(_0371_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5890__A2 (.I(_1127_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5892__A1 (.I(_0500_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5893__A1 (.I(_0578_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5893__A2 (.I(_1096_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5894__A1 (.I(_1136_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5894__A2 (.I(_1170_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5895__A1 (.I(_0614_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5895__A2 (.I(_1060_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5896__I0 (.I(_0570_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5896__S (.I(_1145_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5897__A2 (.I(_1174_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5898__A2 (.I(_1161_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5900__I (.I(\as2650.r123_2[0][5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5901__A1 (.I(_0709_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5901__A2 (.I(_1119_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5903__I (.I(_0683_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5904__A1 (.I(_1180_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5904__A2 (.I(_1146_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5905__A1 (.I(_0690_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5905__A2 (.I(_1146_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5906__A1 (.I(_0718_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5907__A1 (.I(_0505_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5908__A1 (.I(_0670_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5909__A1 (.I(_0698_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5909__A2 (.I(_1096_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5910__A1 (.I(_1136_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5911__A1 (.I(_0668_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5911__A2 (.I(_1060_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5912__I0 (.I(_0662_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5912__S (.I(_1082_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5913__A2 (.I(_1189_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5916__I (.I(\as2650.r123_2[0][6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5917__A1 (.I(_0763_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5918__A1 (.I(_0759_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5918__C (.I(_1165_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5919__A1 (.I(_0753_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5920__A1 (.I(_0639_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5921__A1 (.I(_0751_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5921__B (.I(_1061_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5923__A1 (.I(_0771_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5923__B (.I(_1134_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5924__A1 (.I(_0749_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5924__A2 (.I(_1057_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5924__B (.I(_1145_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5925__A1 (.I(_0740_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5926__A1 (.I(_0781_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5926__A2 (.I(_1119_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5928__A2 (.I(_1201_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5928__C (.I(_1053_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5930__I (.I(\as2650.r123_2[0][7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5931__A1 (.I(_0724_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5931__B (.I(_0794_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5933__B (.I(_0555_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5934__A1 (.I(_0544_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5935__B1 (.I(_0815_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5935__B2 (.I(_0651_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5936__A1 (.I(_0473_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5937__A1 (.I(_0473_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5937__A2 (.I(_0801_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5938__A1 (.I(_0836_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5938__B (.I(_1067_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5939__A1 (.I(_0834_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5939__A2 (.I(_1071_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5940__A1 (.I(_0516_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5940__A2 (.I(_1164_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5941__A1 (.I(_0840_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5941__A2 (.I(_1165_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5941__B (.I(_1215_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5942__A1 (.I(_0680_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5942__A2 (.I(_1127_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5943__A1 (.I(_0789_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5943__A2 (.I(_1110_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5945__A1 (.I(_0830_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5945__A2 (.I(_1059_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5945__B (.I(_1136_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5945__C (.I(_1219_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5946__A1 (.I(_0828_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5946__A2 (.I(_1057_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5948__A1 (.I(_1212_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5949__A1 (.I(_1089_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5949__A2 (.I(_1118_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5950__A2 (.I(_1223_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5950__C (.I(_1053_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5953__A1 (.I(_0876_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5953__A2 (.I(_4157_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5953__A3 (.I(_4278_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5954__I (.I(_1227_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5955__I (.I(_1228_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5957__A1 (.I(_4219_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5957__A2 (.I(_4227_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5958__A1 (.I(_1230_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5958__A2 (.I(_1231_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5959__I (.I(_1232_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5960__I (.I(_4443_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5962__A1 (.I(_4426_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5962__A2 (.I(_1235_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5962__A3 (.I(_4489_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5963__I (.I(_0854_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5964__I (.I(_4197_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5966__A1 (.I(_1238_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5966__A2 (.I(_1239_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5967__A1 (.I(_0469_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5967__A3 (.I(_4432_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5968__I (.I(_4427_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5969__A2 (.I(_1242_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5969__A3 (.I(_4425_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5970__A1 (.I(_1237_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5970__A2 (.I(_1241_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5970__A3 (.I(_1243_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5971__A1 (.I(_1234_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5971__A2 (.I(_1236_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5971__A3 (.I(_1244_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5972__A1 (.I(_1229_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5972__A2 (.I(_1233_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5973__A1 (.I(_0868_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5973__A2 (.I(_4423_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5975__I (.I(_1248_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5976__I (.I(_4417_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5977__I (.I(_1250_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5978__I (.I(_1251_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5979__A1 (.I(_1238_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5980__A1 (.I(\as2650.psl[6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5980__A2 (.I(_4428_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5981__A1 (.I(\as2650.psl[7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5981__A2 (.I(_1239_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5983__A1 (.I(_1253_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5983__A2 (.I(_1256_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5984__A1 (.I(_0814_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5984__A2 (.I(_1252_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5984__A3 (.I(_1257_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5985__A1 (.I(_1249_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5986__I (.I(_4393_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5987__I (.I(_4369_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5988__A1 (.I(_4215_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5988__A2 (.I(_4223_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5989__A2 (.I(_4330_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5991__A1 (.I(_1261_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5991__A2 (.I(_1264_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5991__B (.I(_1233_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5991__C (.I(_1228_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5992__A1 (.I(_1260_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5993__A1 (.I(_4174_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5993__A2 (.I(_4167_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5994__I (.I(_1267_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5995__I (.I(_1236_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5996__A1 (.I(_4201_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5996__A2 (.I(_1268_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5996__A4 (.I(_1237_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5997__I (.I(_4543_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5998__I (.I(_1271_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5999__I (.I(_1243_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6000__A1 (.I(_1272_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6000__A2 (.I(_1273_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6001__I (.I(_0879_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6002__I (.I(_1275_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6003__I (.I(_1276_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6006__A1 (.I(_1278_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6006__A2 (.I(_0418_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6006__A3 (.I(_1279_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6007__A1 (.I(_4430_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6007__A2 (.I(_1280_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6008__A1 (.I(_4214_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6008__A2 (.I(_4250_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6009__I (.I(_1282_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6010__A1 (.I(_1277_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6010__A2 (.I(_1281_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6010__B (.I(_1233_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6010__C (.I(_1283_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6011__A1 (.I(_1270_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6012__A3 (.I(_1266_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6013__I (.I(_1229_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6014__I (.I(_1086_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6015__I (.I(_1288_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6016__A1 (.I(_0670_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6016__A2 (.I(_1289_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6017__I (.I(_0685_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6018__I (.I(_1291_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6019__I (.I(_4443_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6020__I (.I(_1293_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6021__I (.I(_1294_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6022__A1 (.I(_4199_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6022__A2 (.I(_1264_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6023__A1 (.I(_1291_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6024__A2 (.I(_1292_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6024__B (.I(_1295_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6024__C (.I(_1297_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6025__A1 (.I(_1290_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6026__A1 (.I(_1287_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6026__B (.I(_1286_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6027__I (.I(_4438_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6028__I (.I(_1301_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6029__A1 (.I(_1226_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6029__A2 (.I(_1286_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6029__C (.I(_1302_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6033__A1 (.I(_4238_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6033__A3 (.I(_1304_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6033__A4 (.I(_1305_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6034__A2 (.I(_1306_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6035__A1 (.I(_4263_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6037__A1 (.I(_4254_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6037__A2 (.I(_0878_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6038__A3 (.I(_1304_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6038__A4 (.I(_1305_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6039__A1 (.I(_1309_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6039__A2 (.I(_1310_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6039__A3 (.I(_1311_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6040__A1 (.I(_1308_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6040__A2 (.I(_1312_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6041__A1 (.I(_4235_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6041__A2 (.I(_4241_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6042__I (.I(_4232_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6043__I (.I(_1315_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6044__A1 (.I(_1316_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6044__A2 (.I(_1267_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6045__A1 (.I(_1314_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6045__A2 (.I(_1317_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6046__I (.I(_1034_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6047__I (.I(_4214_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6048__A1 (.I(_1320_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6048__A2 (.I(_1228_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6049__I (.I(_1315_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6050__I (.I(_1322_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6051__I (.I(_0889_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6052__A1 (.I(_4174_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6053__A1 (.I(_0883_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6053__A2 (.I(_1325_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6055__A1 (.I(_1316_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6055__A2 (.I(_1327_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6056__I (.I(_4235_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6057__A1 (.I(_1329_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6057__A2 (.I(_1306_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6058__A1 (.I(_1328_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6059__A1 (.I(_1323_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6059__A2 (.I(_1324_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6059__B (.I(_1331_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6060__A1 (.I(_1319_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6060__A2 (.I(_1321_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6061__A1 (.I(_1318_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6061__A2 (.I(_1333_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6062__I (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6063__I (.I(_1335_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6064__A3 (.I(_1304_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6064__A4 (.I(_1305_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6065__A1 (.I(_4238_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6065__A2 (.I(_1337_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6066__A1 (.I(_1336_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6066__A2 (.I(_1338_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6067__I (.I(_0881_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6068__I (.I(_4263_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6069__A1 (.I(_1340_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6070__A1 (.I(_1339_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6070__A2 (.I(_1342_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6070__B (.I(_1323_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6071__A1 (.I(_1322_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6071__A2 (.I(_1086_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6072__A2 (.I(_1344_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6073__I (.I(_4167_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6074__A1 (.I(_1346_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6074__A2 (.I(_4237_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6076__A1 (.I(\as2650.cycle[3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6076__A3 (.I(_4174_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6076__A4 (.I(_4172_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6077__A1 (.I(_0883_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6077__A2 (.I(_1315_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6077__A3 (.I(_1349_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6078__A1 (.I(_1347_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6078__A2 (.I(_1350_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6079__A2 (.I(_1351_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6080__A2 (.I(_1352_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6083__I (.I(_1355_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6084__A1 (.I(_1355_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6084__A2 (.I(_1305_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6085__A1 (.I(_4551_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6085__A2 (.I(_1357_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6086__A1 (.I(_1354_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6086__A2 (.I(_1356_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6086__A3 (.I(_1358_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6087__A1 (.I(_4215_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6088__A2 (.I(_1227_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6089__A1 (.I(_4394_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6089__A2 (.I(_1361_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6090__A1 (.I(_4550_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6090__A2 (.I(_0879_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6091__A1 (.I(_1315_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6091__A2 (.I(_0882_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6092__A1 (.I(_1282_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6092__A2 (.I(_1362_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6092__B (.I(_1363_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6092__C (.I(_1364_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6093__A1 (.I(_1359_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6094__I (.I(_4194_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6095__A1 (.I(_4442_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6095__A2 (.I(_1228_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6096__A1 (.I(_4328_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6096__A2 (.I(_1230_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6098__A1 (.I(_1367_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6098__A2 (.I(_1283_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6098__B1 (.I(_1368_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6098__B2 (.I(_1370_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6099__A2 (.I(_1353_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6099__A3 (.I(_1366_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6099__A4 (.I(_1371_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6100__I (.I(_1372_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6101__I (.I(_1323_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6102__A1 (.I(_1374_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6103__I (.I(_1375_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6104__I (.I(_1375_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6105__A2 (.I(_1100_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6106__A1 (.I(_4441_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6107__I (.I(_1372_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6109__A2 (.I(_1379_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6109__C (.I(_1302_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6110__I (.I(_0337_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6111__I (.I(_4387_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6112__A2 (.I(_1383_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6113__A1 (.I(_1382_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6115__A2 (.I(_1385_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6115__C (.I(_1302_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6116__A2 (.I(_4527_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6117__A1 (.I(_0917_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6119__I (.I(_4202_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6120__I (.I(_1390_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6121__I (.I(_1391_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6122__A2 (.I(_1388_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6122__C (.I(_1392_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6123__I (.I(_0464_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6124__A2 (.I(_1393_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6125__A1 (.I(_0924_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6127__A2 (.I(_1395_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6127__C (.I(_1392_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6128__I (.I(_1372_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6129__I (.I(_1375_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6130__I (.I(_1375_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6131__A1 (.I(_1399_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6131__A2 (.I(_0694_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6132__A1 (.I(_0579_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6133__I (.I(_1372_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6135__A2 (.I(_1401_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6135__C (.I(_1392_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6136__A1 (.I(_1399_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6136__A2 (.I(_0593_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6137__A1 (.I(_0711_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6139__A2 (.I(_1405_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6139__C (.I(_1392_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6140__A1 (.I(_1399_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6140__A2 (.I(_0681_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6141__A1 (.I(_0944_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6143__I (.I(_1391_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6144__A2 (.I(_1408_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6144__C (.I(_1410_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6145__I (.I(_0790_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6146__A1 (.I(_1399_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6146__A2 (.I(_0754_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6147__A1 (.I(_1411_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6148__A1 (.I(net21));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6149__A2 (.I(_1413_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6149__C (.I(_1410_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6150__A1 (.I(_0622_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6150__A2 (.I(_1019_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6152__I (.I(_1416_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6153__I (.I(_1416_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6155__A1 (.I(_0976_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6158__A1 (.I(_0985_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6160__A1 (.I(_0993_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6162__A1 (.I(_1000_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6164__A1 (.I(_1006_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6165__A1 (.I(\as2650.stack[4][13] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6165__A2 (.I(_1416_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6166__A1 (.I(_1012_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6167__A1 (.I(\as2650.stack[4][14] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6167__A2 (.I(_1416_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6168__A1 (.I(_1016_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6169__A1 (.I(_4344_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6169__A2 (.I(_0321_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6169__A3 (.I(_0422_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6169__A4 (.I(_0476_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6170__A1 (.I(_0569_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6170__A2 (.I(_0662_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6170__A3 (.I(_0740_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6171__I (.I(_0548_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6172__A1 (.I(_1429_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6172__A2 (.I(_0753_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6173__A2 (.I(_1429_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6174__A1 (.I(_4303_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6174__A2 (.I(_0403_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6175__A2 (.I(_1432_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6176__A1 (.I(_0442_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6176__A2 (.I(_0467_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6177__A2 (.I(_0561_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6178__A1 (.I(_0641_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6179__A2 (.I(_0795_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6179__A3 (.I(_1436_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6180__A2 (.I(_1431_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6181__A1 (.I(\as2650.psl[1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6181__A2 (.I(_0795_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6182__A1 (.I(_0795_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6184__I (.I(_1234_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6185__I (.I(_1442_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6186__A1 (.I(_4258_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6186__A2 (.I(_1440_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6186__A3 (.I(_1441_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6186__B (.I(_1443_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6187__A1 (.I(_0408_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6187__A3 (.I(_0543_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6187__A4 (.I(_0641_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6188__A1 (.I(_1252_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6188__A2 (.I(_0403_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6188__A3 (.I(_0720_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6188__A4 (.I(_0801_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6189__A1 (.I(_4311_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6189__A2 (.I(_1445_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6190__A2 (.I(_1447_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6191__A1 (.I(_0600_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6191__A2 (.I(_0821_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6191__A3 (.I(_1428_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6192__I (.I(_1374_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6193__I (.I(_1450_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6194__A1 (.I(_1322_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6194__A2 (.I(_0447_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6195__A1 (.I(_0394_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6196__A1 (.I(_0360_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6196__A2 (.I(_4541_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6196__A3 (.I(_4405_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6197__A1 (.I(_0751_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6197__A2 (.I(_0669_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6197__A3 (.I(_0500_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6197__A4 (.I(_0492_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6198__A1 (.I(_1454_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6198__B (.I(_0789_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6199__A1 (.I(_0394_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6200__A1 (.I(_0754_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6200__A2 (.I(_1457_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6201__A1 (.I(_0824_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6202__A1 (.I(_1453_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6202__A2 (.I(_1456_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6202__C (.I(_1295_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6203__A1 (.I(_1451_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6204__I (.I(_4250_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6205__I (.I(_1462_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6206__I (.I(_0884_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6207__A1 (.I(_1464_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6207__A2 (.I(_1355_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6208__A1 (.I(_1320_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6209__A1 (.I(_1465_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6209__A2 (.I(_1232_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6209__A3 (.I(_1466_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6210__A1 (.I(_0393_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6210__A2 (.I(_4431_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6211__A1 (.I(_0340_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6211__A2 (.I(_1468_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6211__B (.I(_1429_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6212__A1 (.I(_4543_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6212__A2 (.I(_1361_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6213__A1 (.I(_4255_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6213__A2 (.I(_4232_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6214__A2 (.I(_4489_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6215__A1 (.I(_1471_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6215__A2 (.I(_0394_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6215__A3 (.I(_1472_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6216__A1 (.I(_1045_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6216__A2 (.I(_1470_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6217__A1 (.I(_1463_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6217__A2 (.I(_1467_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6217__B1 (.I(_1469_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6217__B2 (.I(_1474_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6218__A1 (.I(_1293_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6218__A2 (.I(_0516_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6218__A3 (.I(_1229_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6219__A1 (.I(_1095_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6219__A2 (.I(_1242_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6219__B1 (.I(_4544_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6219__B2 (.I(_4199_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6220__A1 (.I(_4187_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6220__A2 (.I(_1477_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6220__B (.I(_4419_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6221__I (.I(_1465_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6223__A1 (.I(_1320_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6223__A2 (.I(_1250_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6224__I (.I(_0867_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6225__A1 (.I(_1482_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6226__A1 (.I(_1479_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6226__A2 (.I(_4187_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6226__B1 (.I(_1480_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6226__B2 (.I(_1481_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6226__C (.I(_1483_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6227__A1 (.I(_1476_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6227__A3 (.I(_1484_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6228__I (.I(_1034_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6229__A1 (.I(_4551_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6229__A2 (.I(_1271_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6229__A3 (.I(_0397_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6229__A4 (.I(_0339_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6230__A1 (.I(_1486_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6230__A2 (.I(_1487_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6231__I (.I(_0882_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6232__I (.I(_1489_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6233__A1 (.I(_1490_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6233__A2 (.I(_1317_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6234__A2 (.I(_1237_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6235__A1 (.I(_4550_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6235__A2 (.I(_4341_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6235__A3 (.I(_0338_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6235__B (.I(_4417_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6236__A1 (.I(_4544_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6236__A2 (.I(_1453_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6237__A1 (.I(_1323_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6237__A2 (.I(_1493_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6238__A1 (.I(_1316_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6238__A2 (.I(_1275_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6238__B (.I(_1357_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6239__I (.I(_4255_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6240__I (.I(_1497_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6241__A1 (.I(_1498_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6241__A2 (.I(_1248_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6242__I (.I(_4208_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6243__A1 (.I(_0884_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6243__A2 (.I(_4167_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6244__A1 (.I(_1500_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6244__A2 (.I(_1501_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6245__A1 (.I(_4442_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6245__A2 (.I(_1241_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6246__A1 (.I(_0867_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6246__A2 (.I(_4550_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6247__A1 (.I(_1499_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6247__A2 (.I(_1502_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6247__A3 (.I(_1503_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6247__A4 (.I(_1504_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6248__A1 (.I(_1492_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6248__A2 (.I(_1495_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6248__A3 (.I(_1496_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6248__A4 (.I(_1505_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6249__A1 (.I(_1464_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6249__A2 (.I(_0883_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6250__A1 (.I(_1346_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6250__A2 (.I(_1507_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6251__I (.I(_1508_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6252__A1 (.I(_1238_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6253__A1 (.I(_1509_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6253__A2 (.I(_1510_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6254__A1 (.I(_1488_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6254__A2 (.I(_1491_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6255__I (.I(_1471_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6256__A1 (.I(_0814_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6256__A2 (.I(_1513_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6256__A3 (.I(_1266_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6257__A1 (.I(_1475_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6257__A3 (.I(_1512_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6258__I (.I(_1095_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6259__I (.I(_1516_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6260__I (.I(_1517_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6261__I (.I(_1043_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6262__I (.I(_1519_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6263__A1 (.I(_1064_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6263__A2 (.I(_0745_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6264__A1 (.I(_1520_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6264__A2 (.I(_0681_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6265__I (.I(_4428_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6266__I (.I(_1288_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6267__I (.I(\as2650.psl[6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6268__I (.I(_0758_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6269__I (.I(_1280_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6270__A1 (.I(_1239_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6270__A2 (.I(_0759_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6271__A1 (.I(_1525_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6271__A2 (.I(_1526_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6271__B (.I(_1527_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6272__I (.I(_0751_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6273__A1 (.I(_1530_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6273__A2 (.I(_1273_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6274__I (.I(_4418_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6275__A1 (.I(_1273_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6275__A2 (.I(_1456_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6275__C (.I(_1532_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6276__A1 (.I(_1523_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6276__A2 (.I(_1524_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6277__I (.I(_4227_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6278__A1 (.I(_1535_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6278__A2 (.I(_0840_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6279__I (.I(_0718_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6280__A2 (.I(_1537_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6281__A1 (.I(_1383_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6281__A2 (.I(_0754_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6281__A3 (.I(_0481_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6282__A1 (.I(_4328_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6284__A1 (.I(_1045_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6284__A2 (.I(_1534_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6284__B2 (.I(_1539_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6284__C (.I(_1541_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6285__A2 (.I(_1542_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6286__I (.I(_1335_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6287__I (.I(_1544_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6290__A1 (.I(_1546_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6290__A2 (.I(_1547_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6291__I (.I(_4391_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6292__I (.I(_1549_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6293__I (.I(_1550_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6294__I (.I(_4531_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6295__I (.I(_0373_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6296__I (.I(_1553_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6297__I (.I(_1554_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6298__I (.I(_1147_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6299__A1 (.I(_1551_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6299__A2 (.I(_1552_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6299__A3 (.I(_1555_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6299__A4 (.I(_1556_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6300__I (.I(_0597_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6301__I (.I(_1526_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6302__A1 (.I(_1558_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6302__A2 (.I(_1291_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6302__A3 (.I(_1559_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6303__A1 (.I(_1547_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6304__A1 (.I(_1518_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6304__A3 (.I(_1548_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6304__A4 (.I(_1561_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6305__A1 (.I(_1515_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6306__A2 (.I(_1461_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6308__I (.I(_1565_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6309__A1 (.I(_1525_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6309__A2 (.I(_1515_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6309__B (.I(_1566_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6310__A1 (.I(_1564_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6311__A1 (.I(_4258_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6311__A2 (.I(_1212_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6312__I (.I(_1462_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6313__I (.I(_1569_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6314__I (.I(_1532_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6315__I (.I(_1571_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6316__A1 (.I(_1411_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6316__A2 (.I(_1457_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6316__C (.I(_1572_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6317__A1 (.I(_1570_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6318__I (.I(_1374_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6319__I (.I(_1575_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6320__A1 (.I(_1541_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6321__A1 (.I(_1278_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6321__A2 (.I(_4314_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6321__A3 (.I(_1279_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6322__I (.I(_0837_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6323__I (.I(_0595_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6325__I (.I(_1581_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6326__A1 (.I(_4463_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6326__A2 (.I(_1104_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6326__B1 (.I(_0375_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6326__B2 (.I(_0849_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6327__I (.I(net9));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6328__I (.I(_1584_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6330__I (.I(_1586_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6331__I (.I(_1587_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6333__A1 (.I(\as2650.psu[3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6333__A2 (.I(_1585_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6333__B1 (.I(_1588_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6333__B2 (.I(net27));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6333__C1 (.I(_1589_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6333__C2 (.I(_4392_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6334__A1 (.I(_1226_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6334__A2 (.I(_0684_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6335__A1 (.I(\as2650.psu[7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6335__A2 (.I(_1579_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6335__B1 (.I(_1582_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6335__B2 (.I(\as2650.psu[4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6336__A1 (.I(_1523_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6336__A2 (.I(_1578_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6336__A3 (.I(_1592_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6337__I (.I(_1585_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6338__I (.I(\as2650.psl[5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6339__A1 (.I(_4316_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6339__A2 (.I(_4391_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6339__B1 (.I(_0683_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6340__A2 (.I(_0375_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6340__B1 (.I(_1594_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6340__B2 (.I(_4320_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6340__C (.I(_1596_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6341__A1 (.I(\as2650.psl[1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6341__A2 (.I(_1104_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6341__B1 (.I(_1588_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6341__B2 (.I(_1525_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6343__A1 (.I(\as2650.psl[7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6343__A2 (.I(_1599_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6343__B1 (.I(_1581_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6343__B2 (.I(_4248_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6344__I (.I(_1238_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6345__A1 (.I(_1597_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6345__B (.I(_1601_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6346__A1 (.I(_1578_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6346__A2 (.I(_1602_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6347__I (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6348__I (.I(_1604_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6349__A1 (.I(_1549_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6349__A2 (.I(_4334_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6349__B1 (.I(_0592_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6349__B2 (.I(_0684_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6349__C1 (.I(_0753_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6349__C2 (.I(_1605_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6350__A1 (.I(_4530_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6350__A2 (.I(_4387_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6350__B1 (.I(_4526_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6350__B2 (.I(_1554_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6350__C1 (.I(_0680_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6350__C2 (.I(_0758_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6351__A1 (.I(_1147_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6351__A2 (.I(_1393_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6351__B1 (.I(_0505_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6351__B2 (.I(_0597_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6351__C1 (.I(_1578_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6351__C2 (.I(_1601_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6353__A1 (.I(_1261_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6353__A2 (.I(_1527_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6353__B2 (.I(_1609_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6354__I (.I(\as2650.psl[7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6355__I (.I(_1253_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6356__A1 (.I(_1611_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6356__A2 (.I(_1612_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6356__A3 (.I(_1264_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6357__I (.I(_0837_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6358__A1 (.I(_1593_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6358__B2 (.I(_1614_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6359__I (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6361__I (.I(_1617_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6362__I (.I(_1618_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6363__A1 (.I(_1619_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6363__A2 (.I(_1281_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6364__A1 (.I(_1281_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6364__B2 (.I(_1611_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6365__I (.I(_1442_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6366__I (.I(_4219_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6367__I (.I(_1623_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6368__A1 (.I(_1622_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6368__A2 (.I(_1624_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6369__A1 (.I(_0790_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6369__A2 (.I(_1571_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6370__I (.I(_1519_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6371__I (.I(_1480_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6372__A1 (.I(_1520_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6372__A2 (.I(_1537_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6372__B (.I(_1628_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6373__A1 (.I(_1621_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6373__B2 (.I(_1627_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6373__C (.I(_1629_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6375__A1 (.I(_1576_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6375__A2 (.I(_1548_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6376__A2 (.I(_1574_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6377__I (.I(_1565_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6378__I (.I(_1634_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6379__A1 (.I(_1611_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6379__A2 (.I(_1515_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6379__B (.I(_1635_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6380__A1 (.I(_1515_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6380__A2 (.I(_1633_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6381__A2 (.I(_4463_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6382__I (.I(_1637_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6383__I (.I(_1638_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6384__I (.I(_1639_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6385__A2 (.I(_1640_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6385__A3 (.I(_1019_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6390__A1 (.I(_0976_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6390__A2 (.I(_1643_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6393__A1 (.I(_0985_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6393__A2 (.I(_1643_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6395__A1 (.I(_0993_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6395__A2 (.I(_1643_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6397__A1 (.I(_1000_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6397__A2 (.I(_1643_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6399__A1 (.I(_1006_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6400__A1 (.I(\as2650.stack[3][13] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6401__A1 (.I(_1012_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6402__A1 (.I(\as2650.stack[3][14] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6403__A1 (.I(_1016_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6404__I (.I(_0975_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6406__I (.I(_1654_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6408__I (.I(_1656_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6409__A2 (.I(_1657_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6409__A3 (.I(_0960_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6410__I (.I(_1658_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6411__I (.I(_1659_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6412__I (.I(_1659_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6413__A1 (.I(\as2650.stack[2][8] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6413__A2 (.I(_1661_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6414__A1 (.I(_1653_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6415__I (.I(_0984_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6416__I (.I(_1658_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6418__A1 (.I(_1663_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6419__I (.I(_0992_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6420__A1 (.I(\as2650.stack[2][10] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6421__A1 (.I(_1666_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6422__I (.I(_0999_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6423__A1 (.I(\as2650.stack[2][11] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6424__A1 (.I(_1668_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6425__I (.I(_1005_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6426__A1 (.I(\as2650.stack[2][12] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6427__A1 (.I(_1670_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6427__A2 (.I(_1661_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6428__I (.I(_1011_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6429__A1 (.I(\as2650.stack[2][13] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6429__A2 (.I(_1659_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6430__A1 (.I(_1672_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6430__A2 (.I(_1661_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6432__A2 (.I(_1659_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6433__A1 (.I(_1674_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6433__A2 (.I(_1661_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6434__I (.I(_1500_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6435__I (.I(_1676_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6436__I (.I(_1464_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6437__I (.I(_1335_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6438__I (.I(_1679_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6439__A1 (.I(_1253_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6439__A2 (.I(_4431_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6440__A1 (.I(_4223_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6440__A2 (.I(_1681_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6441__A1 (.I(_0876_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6441__A2 (.I(_1682_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6442__I (.I(_1683_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6443__I (.I(_1684_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6444__A1 (.I(_1680_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6444__A2 (.I(_1685_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6445__A1 (.I(_1678_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6446__A1 (.I(_1677_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6446__A2 (.I(_1118_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6446__A3 (.I(_1356_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6446__A4 (.I(_1687_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6447__I (.I(_1688_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6449__I (.I(_1551_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6450__I (.I(_1502_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6451__A1 (.I(_1691_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6451__A2 (.I(_1692_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6451__B (.I(_1690_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6452__A1 (.I(_1523_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6452__A2 (.I(_1690_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6453__A1 (.I(_1552_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6453__A2 (.I(_1692_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6454__A1 (.I(_1239_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6454__A2 (.I(_1690_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6455__I (.I(_0877_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6457__A1 (.I(_1678_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6457__A2 (.I(_1354_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6457__A3 (.I(_0852_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6457__A4 (.I(_1346_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6458__I (.I(_1697_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6459__I (.I(_1554_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6460__A1 (.I(_1696_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6460__A2 (.I(_1688_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6460__B1 (.I(_1698_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6460__B2 (.I(_1699_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6462__I (.I(_1504_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6463__A1 (.I(_1502_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6463__A2 (.I(_1701_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6464__A1 (.I(_1292_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6464__A2 (.I(_1692_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6464__B (.I(_1702_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6465__I (.I(_1697_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6466__A1 (.I(_0814_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6466__A2 (.I(_1704_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6467__A1 (.I(_1690_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6468__I (.I(_1559_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6469__A1 (.I(_4160_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6469__A2 (.I(_1688_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6469__B1 (.I(_1698_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6469__B2 (.I(_1706_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6471__I (.I(_1604_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6472__I (.I(_1708_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6473__I (.I(_1709_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6474__I (.I(_1710_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6475__A1 (.I(_4328_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6475__A2 (.I(_1688_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6475__B1 (.I(_1704_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6475__B2 (.I(_1711_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6476__I (.I(_1712_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6477__I (.I(_1084_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6478__A1 (.I(_1601_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6478__A2 (.I(_1051_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6480__A1 (.I(_0853_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6480__A2 (.I(_4489_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6482__A1 (.I(_1716_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6482__A2 (.I(_1035_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6482__B (.I(_1717_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6482__C (.I(_4202_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6484__I0 (.I(\as2650.r123[0][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6484__I1 (.I(\as2650.r123_2[0][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6485__I (.I(_1720_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6486__I (.I(_1721_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6488__A1 (.I(_4405_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6489__A1 (.I(_0294_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6489__A2 (.I(_4152_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6489__A3 (.I(_4419_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6489__A4 (.I(_1236_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6492__A2 (.I(_1719_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6492__B2 (.I(_1727_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6493__A2 (.I(_1715_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6495__I0 (.I(\as2650.r123[0][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6495__I1 (.I(\as2650.r123_2[0][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6496__I (.I(_1730_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6498__I (.I(_1732_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6499__A1 (.I(_4541_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6499__A2 (.I(_1733_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6502__A1 (.I(_0337_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6502__A2 (.I(_1736_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6502__B1 (.I(_1733_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6502__B2 (.I(_4441_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6503__A1 (.I(_1735_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6504__A1 (.I(\as2650.r123_2[1][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6504__A2 (.I(_1729_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6504__B1 (.I(_1727_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6504__B2 (.I(_1738_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6505__A1 (.I(_1116_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6505__A2 (.I(_1717_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6508__A1 (.I(_0359_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6509__A1 (.I(_4541_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6509__A2 (.I(_1733_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6510__I0 (.I(\as2650.r123[0][2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6510__I1 (.I(\as2650.r123_2[0][2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6511__I (.I(_1744_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6512__I (.I(_1745_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6513__A1 (.I(_4284_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6514__I (.I(_1745_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6516__A1 (.I(_4383_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6516__A3 (.I(_1732_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6516__A4 (.I(_1749_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6520__A2 (.I(_1719_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6520__B1 (.I(_1741_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6520__B2 (.I(_1753_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6521__A1 (.I(_1139_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6521__A2 (.I(_1715_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6522__A1 (.I(_0364_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6525__A1 (.I(_1757_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6526__I (.I(\as2650.r0[2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6527__A1 (.I(_1759_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6528__I0 (.I(\as2650.r123[0][3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6528__I1 (.I(\as2650.r123_2[0][3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6528__S (.I(_4144_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6529__I (.I(_1761_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6531__I (.I(_1763_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6532__A1 (.I(_4405_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6532__A2 (.I(_1764_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6535__A1 (.I(_0359_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6540__A2 (.I(_1719_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6540__B1 (.I(_1741_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6540__B2 (.I(_1772_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6541__A1 (.I(_1156_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6541__A2 (.I(_1715_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6544__A1 (.I(_1757_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6544__A2 (.I(_1763_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6545__A1 (.I(_0363_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6545__A2 (.I(_1732_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6546__A1 (.I(_1759_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6546__A2 (.I(_1749_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6548__A2 (.I(\as2650.r123_2[0][4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6549__A1 (.I(_4147_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6549__A2 (.I(_0540_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6550__A1 (.I(_4285_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6550__A2 (.I(_1781_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6552__A1 (.I(_4382_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6552__B2 (.I(_4284_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6553__B1 (.I(_1784_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6554__A1 (.I(_0499_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6554__A2 (.I(_1721_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6555__A2 (.I(_1785_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6556__A1 (.I(_0492_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6558__A1 (.I(_1779_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6561__A2 (.I(_1719_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6561__B1 (.I(_1741_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6562__A1 (.I(_1174_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6562__A2 (.I(_1715_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6564__I (.I(_1794_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6568__A1 (.I(_1779_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6570__A1 (.I(_1779_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6571__A1 (.I(_1785_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6572__A1 (.I(_1785_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6574__A1 (.I(_4519_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6575__A1 (.I(_0498_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6576__A1 (.I(_0363_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6577__A3 (.I(_1807_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6578__I0 (.I(\as2650.r123[0][5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6578__I1 (.I(\as2650.r123_2[0][5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6578__S (.I(_4144_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6579__I (.I(_1809_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6581__I (.I(_1811_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6582__A2 (.I(_1812_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6584__A1 (.I(_4383_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6584__A2 (.I(_1781_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6585__A1 (.I(_1759_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6585__B2 (.I(_1757_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6587__A1 (.I(_0585_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6587__A2 (.I(_1721_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6593__A1 (.I(_1795_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6593__A2 (.I(_1823_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6594__A2 (.I(_1729_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6595__A1 (.I(_1189_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6598__A1 (.I(_1785_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6604__A1 (.I(_0669_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6604__A2 (.I(_1736_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6605__A1 (.I(_0669_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6608__A2 (.I(_1812_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6609__A1 (.I(_4382_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6609__A2 (.I(_1811_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6610__I0 (.I(\as2650.r123[0][6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6610__I1 (.I(\as2650.r123_2[0][6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6611__I (.I(_1840_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6612__A1 (.I(\as2650.r0[0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6613__A1 (.I(_4382_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6613__A2 (.I(_4284_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6615__A1 (.I(\as2650.r0[3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6616__A1 (.I(\as2650.r0[5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6616__A2 (.I(_1730_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6617__A1 (.I(\as2650.r0[4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6617__A2 (.I(_1745_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6618__A1 (.I(_1845_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6619__A1 (.I(_1844_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6620__A1 (.I(_4520_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6620__A2 (.I(_1781_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6621__A1 (.I(_0363_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6621__B1 (.I(_1763_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6621__B2 (.I(_1759_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6622__A2 (.I(_1845_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6623__A1 (.I(_0671_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6623__A2 (.I(_1721_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6626__A2 (.I(_1849_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6629__A3 (.I(_1858_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6630__A1 (.I(_1795_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6630__A2 (.I(_1859_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6631__A2 (.I(_1729_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6632__A1 (.I(_1201_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6632__A2 (.I(_1717_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6634__A2 (.I(_1858_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6635__A2 (.I(_1858_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6642__A2 (.I(_1849_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6643__A2 (.I(_1849_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6645__A1 (.I(_1844_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6646__A1 (.I(_0671_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6647__A1 (.I(\as2650.r0[4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6648__A1 (.I(\as2650.r0[5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6648__A2 (.I(_1745_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6651__A2 (.I(_1840_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6652__A1 (.I(\as2650.r0[2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6652__A2 (.I(_1809_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6653__I0 (.I(\as2650.r123[0][7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6653__I1 (.I(\as2650.r123_2[0][7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6653__S (.I(_4144_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6654__A1 (.I(\as2650.r0[0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6654__A2 (.I(_1882_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6657__A2 (.I(_1879_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6657__A3 (.I(_1885_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6658__I (.I(_1781_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6659__A1 (.I(_0364_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6659__A2 (.I(_1887_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6660__A1 (.I(_0498_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6660__B2 (.I(_0362_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6661__A1 (.I(_1807_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6662__A2 (.I(_1720_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6668__A2 (.I(_1896_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6670__A1 (.I(_1795_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6670__A2 (.I(_1898_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6671__A2 (.I(_1729_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6672__A1 (.I(_1223_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6672__A2 (.I(_1717_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6675__I (.I(_1902_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6677__I (.I(_1904_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6678__A1 (.I(_0866_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6678__A2 (.I(_1905_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6678__A3 (.I(_0960_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6680__I (.I(_1907_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6681__I (.I(_1907_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6682__A2 (.I(_1909_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6683__A1 (.I(_1653_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6683__A2 (.I(_1908_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6686__A1 (.I(_1663_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6686__A2 (.I(_1908_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6688__A1 (.I(_1666_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6688__A2 (.I(_1908_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6690__A1 (.I(_1668_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6690__A2 (.I(_1908_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6691__A1 (.I(\as2650.stack[1][12] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6692__A1 (.I(_1670_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6692__A2 (.I(_1909_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6693__A2 (.I(_1907_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6694__A1 (.I(_1672_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6694__A2 (.I(_1909_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6695__A2 (.I(_1907_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6696__A1 (.I(_1674_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6696__A2 (.I(_1909_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6697__A2 (.I(_4458_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6698__I (.I(_1918_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6699__I (.I(_1919_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6700__I (.I(_1920_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6701__A1 (.I(_0866_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6701__A2 (.I(_1921_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6701__A3 (.I(_0960_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6702__I (.I(_1922_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6703__I (.I(_1923_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6704__I (.I(_1923_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6706__A1 (.I(_1653_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6707__I (.I(_1922_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6708__A1 (.I(\as2650.stack[0][9] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6709__A1 (.I(_1663_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6710__A1 (.I(\as2650.stack[0][10] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6711__A1 (.I(_1666_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6712__A1 (.I(\as2650.stack[0][11] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6713__A1 (.I(_1668_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6714__A1 (.I(\as2650.stack[0][12] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6715__A1 (.I(_1670_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6716__A2 (.I(_1923_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6717__A1 (.I(_1672_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6718__A2 (.I(_1923_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6719__A1 (.I(_1674_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6720__A1 (.I(_1059_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6720__A2 (.I(_1145_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6720__A3 (.I(_1165_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6721__A1 (.I(_4195_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6721__A2 (.I(_1164_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6722__A2 (.I(_1215_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6723__A1 (.I(_1934_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6723__B (.I(_1261_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6725__I (.I(_1716_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6726__A1 (.I(_1612_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6726__A2 (.I(_1051_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6727__A1 (.I(_1939_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6727__A2 (.I(_1035_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6727__B (.I(_1940_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6727__C (.I(_4438_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6729__A2 (.I(_1896_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6734__A1 (.I(_0788_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6734__A2 (.I(_1736_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6736__A1 (.I(_1879_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6736__A2 (.I(_1885_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6737__A1 (.I(_1879_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6737__A2 (.I(_1885_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6739__A1 (.I(\as2650.r0[5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6739__A2 (.I(_1761_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6741__A1 (.I(_0672_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6741__A2 (.I(_1732_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6743__A1 (.I(_0499_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6743__A2 (.I(_1887_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6746__A1 (.I(_1879_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6746__A2 (.I(_1885_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6747__A2 (.I(_1730_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6748__A1 (.I(\as2650.r0[6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6748__A2 (.I(_1744_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6751__I (.I(_1882_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6755__A1 (.I(\as2650.r0[3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6756__I (.I(_1840_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6757__A1 (.I(_4519_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6763__A1 (.I(_1949_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6765__A1 (.I(_1944_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6766__I (.I(_1741_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6767__A2 (.I(_1942_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6767__B1 (.I(_1979_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6767__B2 (.I(_1980_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6768__A2 (.I(_1938_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6769__A1 (.I(_1116_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6769__A2 (.I(_1940_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6769__B1 (.I(_1942_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6771__A1 (.I(_1944_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6773__A1 (.I(_1949_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6780__A1 (.I(_0586_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6780__A2 (.I(_1887_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6787__A2 (.I(_1749_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6787__B1 (.I(_1764_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6787__B2 (.I(_0672_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6788__A2 (.I(_1763_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6789__A2 (.I(_2001_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6791__A1 (.I(_4519_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6793__A1 (.I(_1757_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6793__B2 (.I(_4520_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6795__A1 (.I(_0362_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6796__A1 (.I(_0498_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6796__A2 (.I(_1811_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6805__A1 (.I(_1727_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6805__A2 (.I(_2017_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6815__I (.I(_1887_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6816__A1 (.I(_2027_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6817__A1 (.I(_0750_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6817__A2 (.I(_2027_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6823__A1 (.I(_0362_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6826__A1 (.I(\as2650.r0[4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6827__A1 (.I(_0585_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6830__A1 (.I(_2001_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6836__A1 (.I(_2021_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6837__A2 (.I(_2019_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6837__B2 (.I(_1980_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6838__A1 (.I(_1139_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6838__A2 (.I(_1938_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6840__A1 (.I(_2021_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6847__A1 (.I(_0788_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6847__A2 (.I(_2027_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6848__A1 (.I(_0499_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6849__A1 (.I(_0671_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6849__A2 (.I(_1811_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6850__A1 (.I(_0585_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6856__A1 (.I(_4367_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6856__A2 (.I(_1764_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6866__A2 (.I(_2019_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6866__B1 (.I(_2076_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6866__B2 (.I(_1980_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6867__A1 (.I(_1156_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6867__A2 (.I(_1938_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6873__A1 (.I(_0586_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6875__A1 (.I(_0750_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6875__A2 (.I(_2084_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6877__A1 (.I(_4367_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6877__A2 (.I(_1812_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6888__A1 (.I(_2021_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6891__A1 (.I(_1794_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6891__A2 (.I(_2100_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6892__A2 (.I(_1942_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6893__A1 (.I(_1174_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6893__A2 (.I(_1938_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6901__A1 (.I(_0750_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6901__A2 (.I(_2109_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6903__A1 (.I(_0788_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6903__A2 (.I(_2084_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6906__A2 (.I(_2114_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6909__A2 (.I(_2019_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6909__B2 (.I(_1980_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6910__A1 (.I(_1189_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6911__A1 (.I(_1201_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6911__A2 (.I(_1940_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6911__B1 (.I(_1942_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6915__A2 (.I(_2114_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6916__A1 (.I(_0789_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6916__A2 (.I(_2109_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6918__A2 (.I(_2114_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6922__A1 (.I(_1727_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6922__A2 (.I(_2129_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6924__A2 (.I(_2114_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6926__A1 (.I(_0791_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6926__A2 (.I(_2109_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6927__A1 (.I(_0752_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6927__A2 (.I(_2084_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6930__A1 (.I(_1223_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6930__A2 (.I(_1940_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6930__B1 (.I(_2019_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6931__A1 (.I(_1795_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6932__I (.I(_4295_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6933__I (.I(_0850_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6934__A2 (.I(_1640_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6935__A1 (.I(_0967_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6936__I (.I(_2141_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6938__I (.I(_0862_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6940__I (.I(_2145_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6941__I (.I(_2146_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6942__I (.I(_0957_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6943__I (.I(_0873_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6944__I (.I(_0868_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6945__A1 (.I(_2150_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6945__A2 (.I(_4176_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6946__A1 (.I(_1335_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6947__I (.I(_0881_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6948__I (.I(_0895_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6949__A1 (.I(_1500_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6949__A2 (.I(_1309_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6949__B (.I(_2154_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6950__A1 (.I(_0868_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6950__A2 (.I(_1682_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6951__I (.I(_2156_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6952__A1 (.I(_2153_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6952__A2 (.I(_0889_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6952__B (.I(_2155_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6952__C (.I(_2157_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6953__A1 (.I(_2152_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6954__I (.I(_0898_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6955__A1 (.I(_2149_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6955__A2 (.I(_0875_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6955__A3 (.I(_2159_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6955__B1 (.I(_0897_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6955__B2 (.I(_2160_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6956__A2 (.I(_2161_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6957__A2 (.I(_1657_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6957__A3 (.I(_2162_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6958__I (.I(_2163_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6959__I (.I(_0900_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6960__A2 (.I(_1657_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6962__I (.I(_2167_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6963__A1 (.I(_2147_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6963__B2 (.I(\as2650.stack[2][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6964__A1 (.I(_2138_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6965__I (.I(_0912_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6966__I (.I(_2163_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6967__I (.I(_2167_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6968__I (.I(_2141_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6969__A1 (.I(_2170_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6969__A2 (.I(_2171_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6969__C (.I(_2173_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6970__I (.I(_0858_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6972__A1 (.I(_0908_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6972__A2 (.I(_2176_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6975__A1 (.I(_2178_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6975__A2 (.I(_2171_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6975__C (.I(_2173_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6976__A1 (.I(_0918_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6976__A2 (.I(_2176_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6979__I (.I(_2181_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6980__I (.I(_2182_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6981__A1 (.I(_2183_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6981__A2 (.I(_2171_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6981__C (.I(_2173_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6982__A1 (.I(_0925_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6982__A2 (.I(_2176_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6984__I (.I(_0617_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6986__I (.I(_2187_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6987__I (.I(_2188_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6989__I (.I(_2190_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6990__A1 (.I(_2191_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6991__A1 (.I(_2186_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6994__I (.I(_2194_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6996__I (.I(_2196_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6997__A1 (.I(_2197_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6998__A1 (.I(_2193_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6999__I (.I(_1530_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7000__I (.I(_2199_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7001__I (.I(_0947_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7002__A1 (.I(_2201_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7002__C (.I(_2173_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7003__A1 (.I(_2200_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7004__I (.I(\as2650.pc[7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7005__I (.I(_2203_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7006__I (.I(_2204_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7007__A1 (.I(_2205_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7007__A2 (.I(_2171_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7007__C (.I(_2141_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7008__A1 (.I(_0951_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7008__A2 (.I(_2176_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7010__A1 (.I(_1118_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7010__A2 (.I(_1009_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7011__A2 (.I(_2208_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7012__I (.I(_2209_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7014__I (.I(_2162_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7015__A1 (.I(_0622_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7016__I (.I(_2213_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7017__I (.I(_4474_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7018__A1 (.I(_2215_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7018__A2 (.I(_0901_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7019__I (.I(_2216_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7020__A1 (.I(_2147_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7020__B1 (.I(_2217_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7020__B2 (.I(\as2650.stack[4][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7021__A1 (.I(_2138_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7022__I (.I(_2213_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7023__I (.I(_2216_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7024__I (.I(_2209_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7025__A1 (.I(_2170_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7025__A2 (.I(_2219_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7025__B1 (.I(_2220_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7025__C (.I(_2221_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7026__I (.I(_0957_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7027__A1 (.I(_2223_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7027__A2 (.I(_4482_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7027__A3 (.I(_0968_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7028__A1 (.I(_0908_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7028__A2 (.I(_2224_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7030__A1 (.I(_2178_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7030__A2 (.I(_2219_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7030__B1 (.I(_2220_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7030__B2 (.I(\as2650.stack[4][2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7030__C (.I(_2221_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7031__A1 (.I(_0918_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7031__A2 (.I(_2224_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7033__A1 (.I(_2183_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7033__A2 (.I(_2219_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7033__B1 (.I(_2220_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7033__C (.I(_2221_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7034__A1 (.I(_0925_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7034__A2 (.I(_2224_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7036__A1 (.I(_2191_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7036__B1 (.I(_2217_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7037__A1 (.I(_2186_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7038__A1 (.I(_2197_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7038__B1 (.I(_2217_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7039__A1 (.I(_2193_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7040__A1 (.I(_2201_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7040__B1 (.I(_2217_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7040__B2 (.I(\as2650.stack[4][6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7040__C (.I(_2221_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7041__A1 (.I(_2200_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7042__A1 (.I(_2205_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7042__A2 (.I(_2219_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7042__B1 (.I(_2220_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7042__C (.I(_2209_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7043__A1 (.I(_0951_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7043__A2 (.I(_2224_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7061__A1 (.I(_0967_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7062__I (.I(_2243_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7064__A2 (.I(_1905_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7064__A3 (.I(_2162_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7065__I (.I(_2246_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7066__A2 (.I(_1905_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7067__A2 (.I(_2248_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7068__I (.I(_2249_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7069__A1 (.I(_2147_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7069__B2 (.I(\as2650.stack[1][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7070__A1 (.I(_2138_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7071__I (.I(_2246_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7072__I (.I(_2249_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7073__I (.I(_2243_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7074__A1 (.I(_2170_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7074__B2 (.I(\as2650.stack[1][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7074__C (.I(_2254_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7076__A1 (.I(_0908_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7076__A2 (.I(_2256_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7078__I (.I(_0921_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7079__A1 (.I(_2258_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7079__B2 (.I(\as2650.stack[1][2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7079__C (.I(_2254_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7080__A1 (.I(_0918_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7080__A2 (.I(_2256_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7082__A1 (.I(_2183_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7082__C (.I(_2254_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7083__A1 (.I(_0925_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7083__A2 (.I(_2256_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7085__A1 (.I(_2191_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7086__A1 (.I(_2186_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7087__A1 (.I(_2197_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7087__B2 (.I(\as2650.stack[1][5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7088__A1 (.I(_2193_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7089__I (.I(_0947_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7090__A1 (.I(_2265_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7090__C (.I(_2254_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7091__A1 (.I(_2200_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7092__A1 (.I(_2205_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7092__B2 (.I(\as2650.stack[1][7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7092__C (.I(_2243_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7093__A1 (.I(_0951_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7093__A2 (.I(_2256_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7111__A1 (.I(_0622_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7111__A2 (.I(_2208_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7112__I (.I(_2277_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7114__A2 (.I(_1640_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7115__I (.I(_2280_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7117__I (.I(_2282_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7118__A1 (.I(_2147_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7118__B2 (.I(\as2650.stack[3][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7119__A1 (.I(_2138_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7120__I (.I(_0912_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7121__I (.I(_2280_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7122__I (.I(_2282_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7123__I (.I(_2277_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7124__A1 (.I(_2285_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7124__A2 (.I(_2286_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7124__C (.I(_2288_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7125__I (.I(_1382_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7126__A1 (.I(_2215_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7127__A1 (.I(_2290_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7127__A2 (.I(_2291_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7129__A1 (.I(_2258_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7129__A2 (.I(_2286_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7129__C (.I(_2288_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7130__I (.I(_0917_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7131__A1 (.I(_2294_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7131__A2 (.I(_2291_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7133__I (.I(_2182_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7134__A1 (.I(_2296_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7134__A2 (.I(_2286_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7134__B2 (.I(\as2650.stack[3][3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7134__C (.I(_2288_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7135__I (.I(_0924_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7136__A1 (.I(_2298_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7136__A2 (.I(_2291_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7138__I (.I(_2190_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7139__A1 (.I(_2300_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7139__B2 (.I(\as2650.stack[3][4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7140__A1 (.I(_2186_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7141__I (.I(_2196_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7142__A1 (.I(_2302_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7142__B2 (.I(\as2650.stack[3][5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7143__A1 (.I(_2193_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7144__A1 (.I(_2265_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7144__C (.I(_2288_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7145__A1 (.I(_2200_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7146__I (.I(_2204_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7147__A1 (.I(_2305_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7147__A2 (.I(_2286_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7147__B2 (.I(\as2650.stack[3][7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7147__C (.I(_2277_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7148__I (.I(_1411_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7149__A1 (.I(_2307_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7149__A2 (.I(_2291_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7151__A2 (.I(_2248_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7152__I (.I(_2309_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7154__A2 (.I(_1921_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7154__A3 (.I(_2162_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7155__I (.I(_2312_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7156__A2 (.I(_1921_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7158__I (.I(_2315_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7159__A1 (.I(_2146_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7160__A1 (.I(_0848_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7161__I (.I(_2312_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7162__I (.I(_2315_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7163__I (.I(_2309_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7164__A1 (.I(_2285_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7164__C (.I(_2320_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7165__A2 (.I(_2248_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7166__A1 (.I(_2290_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7168__A1 (.I(_2258_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7168__C (.I(_2320_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7169__A1 (.I(_2294_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7171__A1 (.I(_2296_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7171__B2 (.I(\as2650.stack[0][3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7171__C (.I(_2320_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7172__A1 (.I(_2298_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7174__A1 (.I(_2300_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7175__A1 (.I(_0932_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7176__A1 (.I(_2302_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7177__A1 (.I(_0938_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7178__A1 (.I(_2265_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7178__C (.I(_2320_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7179__A1 (.I(_2199_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7180__A1 (.I(_2305_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7180__C (.I(_2309_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7181__A1 (.I(_2307_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7185__I (.I(_1272_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7187__A1 (.I(_2336_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7187__A2 (.I(_4241_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7188__I (.I(_2337_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7189__A1 (.I(_2335_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7189__A2 (.I(_2338_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7189__A3 (.I(_1324_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7190__I (.I(_1338_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7191__A1 (.I(_1317_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7191__A2 (.I(_2340_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7191__B (.I(_1496_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7192__A1 (.I(_2150_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7192__A2 (.I(_1532_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7192__B (.I(_0871_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7193__A1 (.I(_0852_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7193__A2 (.I(_1283_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7193__A3 (.I(_4253_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7194__A1 (.I(_1351_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7194__A2 (.I(_2341_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7194__A3 (.I(_2342_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7195__A1 (.I(_1086_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7195__A2 (.I(_1683_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7196__A1 (.I(_1500_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7196__A2 (.I(_1349_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7197__A1 (.I(_4393_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7197__A2 (.I(_2156_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7199__A1 (.I(_1464_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7199__A2 (.I(_2348_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7200__A1 (.I(_2156_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7200__A2 (.I(_1310_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7200__A3 (.I(_2346_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7200__B2 (.I(_2349_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7201__A1 (.I(_2345_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7202__A1 (.I(_0877_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7202__A2 (.I(_1260_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7203__I (.I(_2352_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7204__I (.I(_1682_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7205__A1 (.I(_1524_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7205__A2 (.I(_2353_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7205__B (.I(_2354_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7206__A1 (.I(_2351_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7206__B (.I(_1701_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7207__A1 (.I(_1569_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7207__C (.I(_2356_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7208__I (.I(_2357_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7209__I (.I(_2357_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7210__A1 (.I(_1691_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7211__A1 (.I(_2334_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7211__A2 (.I(_2358_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7211__B (.I(_2360_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7212__I (.I(\as2650.addr_buff[1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7213__I (.I(_2361_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7214__I (.I(_2357_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7215__A1 (.I(_2362_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7215__A2 (.I(_2363_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7216__A1 (.I(_1104_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7216__A2 (.I(_2358_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7218__I (.I(_2365_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7219__A1 (.I(_2366_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7219__A2 (.I(_2363_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7220__A1 (.I(_0376_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7220__A2 (.I(_2358_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7221__I (.I(\as2650.addr_buff[3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7222__I (.I(_2368_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7223__I (.I(_2357_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7224__A1 (.I(_1556_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7225__A1 (.I(_2369_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7225__A2 (.I(_2370_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7226__I (.I(\as2650.addr_buff[4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7227__I (.I(_1558_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7228__A1 (.I(_2373_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7229__A1 (.I(_2372_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7229__A2 (.I(_2370_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7230__A1 (.I(_1292_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7231__A2 (.I(_2370_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7232__A1 (.I(_1706_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7232__A2 (.I(_2363_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7233__A1 (.I(_4357_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7233__A2 (.I(_2370_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7234__I (.I(_1579_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7235__A1 (.I(_1340_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7235__A2 (.I(_2363_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7236__A1 (.I(_2377_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7236__A2 (.I(_2358_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7237__A1 (.I(_1309_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7237__A2 (.I(_1491_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7238__A1 (.I(_4179_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7239__A1 (.I(_1252_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7239__A2 (.I(_2380_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7240__I (.I(_1479_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7241__I (.I(_2382_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7242__I (.I(_1489_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7244__I (.I(_2385_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7245__I (.I(_1466_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7246__I (.I(_2387_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7247__A1 (.I(_2383_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7247__A2 (.I(_2386_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7247__A3 (.I(_2380_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7247__A4 (.I(_2388_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7248__A1 (.I(_1367_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7248__A2 (.I(_1279_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7248__A3 (.I(_2346_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7249__I (.I(_1321_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7250__A1 (.I(_1486_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7250__A2 (.I(_2391_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7250__A3 (.I(_1702_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7251__A1 (.I(_2381_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7251__A2 (.I(_2389_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7251__A3 (.I(_2390_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7252__A1 (.I(_1366_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7252__A2 (.I(_2379_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7252__A3 (.I(_2393_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7253__I (.I(_4176_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7254__I (.I(_2395_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7255__A1 (.I(_1451_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7255__A2 (.I(_2396_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7255__B (.I(_1350_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7256__A1 (.I(net24));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7257__A2 (.I(_2397_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7257__C (.I(_1410_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7258__I (.I(_1571_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7259__A1 (.I(_1319_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7259__A2 (.I(_1347_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7260__A1 (.I(_2399_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7260__A2 (.I(_1278_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7260__A3 (.I(_1242_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7260__A4 (.I(_2400_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7261__A2 (.I(_2401_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7262__A1 (.I(_4323_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7262__A2 (.I(_2401_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7262__C (.I(_1410_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7263__I (.I(_1327_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7264__A1 (.I(_1282_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7264__A2 (.I(_1361_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7265__A1 (.I(_2383_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7265__A2 (.I(_1547_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7266__I (.I(_1325_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7267__I (.I(_2406_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7268__I (.I(_1321_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7269__A1 (.I(_1260_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7269__A2 (.I(_1248_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7270__I (.I(_0896_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7271__A1 (.I(_1356_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7271__A2 (.I(_1513_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7271__A3 (.I(_2410_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7271__A4 (.I(_1370_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7272__A1 (.I(_2407_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7272__A2 (.I(_2408_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7272__B1 (.I(_1483_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7272__C (.I(_2411_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7273__A1 (.I(_2403_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7273__B (.I(_2412_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7273__C (.I(_2400_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7274__A1 (.I(net23));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7274__A2 (.I(_2413_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7275__A2 (.I(_2413_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7275__C (.I(_1566_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7276__I (.I(_1301_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7277__I (.I(_2415_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7279__I (.I(_2417_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7280__A1 (.I(_4199_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7280__A2 (.I(_4544_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7281__A1 (.I(_0654_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7281__A2 (.I(_1493_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7281__A3 (.I(_2419_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7282__A1 (.I(_4551_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7282__A2 (.I(_1501_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7283__A1 (.I(_2420_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7284__A1 (.I(_4427_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7284__A3 (.I(_4425_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7285__A1 (.I(_0654_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7285__A2 (.I(_1253_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7285__A3 (.I(_1468_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7285__B (.I(_2423_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7286__A1 (.I(_2419_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7286__A2 (.I(_2424_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7286__B (.I(_4418_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7287__A1 (.I(_2422_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7287__A2 (.I(_2425_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7288__A1 (.I(_1471_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7288__A2 (.I(_1501_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7289__A1 (.I(_1230_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7289__A2 (.I(_2427_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7289__B (.I(_1350_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7290__A1 (.I(_1095_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7290__A2 (.I(_1324_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7291__A1 (.I(_1939_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7291__A3 (.I(_1347_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7292__A1 (.I(_1163_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7292__A2 (.I(_2408_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7292__B (.I(_2406_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7293__A2 (.I(_4237_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7294__A1 (.I(_1355_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7295__A1 (.I(_1312_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7295__A2 (.I(_2433_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7296__A1 (.I(_4233_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7297__A1 (.I(_1314_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7297__A2 (.I(_2435_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7298__A1 (.I(_1497_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7298__A2 (.I(_4543_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7299__I (.I(_0869_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7300__A1 (.I(_4423_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7300__A2 (.I(_1257_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7301__A1 (.I(_4431_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7301__A2 (.I(_1256_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7301__B (.I(_2439_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7302__A2 (.I(_2438_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7302__A3 (.I(_2440_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7303__A1 (.I(_4200_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7303__A2 (.I(_1364_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7303__A3 (.I(_1363_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7304__A1 (.I(_1497_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7304__A2 (.I(_4250_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7305__A1 (.I(_1346_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7305__A2 (.I(_1683_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7305__A3 (.I(_2443_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7306__A1 (.I(_2436_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7306__A2 (.I(_2441_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7306__A3 (.I(_2442_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7306__A4 (.I(_2444_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7307__A1 (.I(_4422_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7307__A2 (.I(_4430_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7307__A3 (.I(_4432_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7307__A4 (.I(_1470_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7308__A1 (.I(_1087_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7308__A2 (.I(_2446_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7309__A1 (.I(_1230_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7309__A2 (.I(_1471_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7309__A3 (.I(_1231_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7309__A4 (.I(_1368_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7310__A1 (.I(_0469_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7310__A2 (.I(_1261_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7310__A3 (.I(_4425_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7311__A1 (.I(_4442_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7311__A2 (.I(_2449_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7312__A1 (.I(_4220_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7312__A2 (.I(_2406_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7312__B (.I(_0970_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7313__A1 (.I(_2450_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7313__A2 (.I(_1503_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7313__A3 (.I(_2451_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7314__A1 (.I(_2406_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7314__A2 (.I(_2448_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7315__A1 (.I(_1501_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7315__A2 (.I(_1504_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7315__A3 (.I(_2351_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7315__B (.I(_2453_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7316__A1 (.I(_2445_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7317__A1 (.I(_2428_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7317__A2 (.I(_2430_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7318__A1 (.I(_1316_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7318__A2 (.I(_4443_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7318__A3 (.I(_0397_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7318__A4 (.I(_0339_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7320__A1 (.I(_4398_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7320__A2 (.I(_1106_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7320__A3 (.I(_0378_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7321__A1 (.I(_0512_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7321__A2 (.I(_0603_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7321__A3 (.I(_0690_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7322__A1 (.I(_4161_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7322__A2 (.I(_2458_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7322__A3 (.I(_0833_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7323__A2 (.I(_2438_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7323__A3 (.I(_2461_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7325__A2 (.I(_2456_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7325__A3 (.I(_2463_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7326__I (.I(_2464_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7327__I (.I(_2465_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7328__I (.I(_1308_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7331__A1 (.I(_2469_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7331__A2 (.I(_4352_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7332__A1 (.I(_1550_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7334__I (.I(_2472_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7335__A2 (.I(_4361_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7336__A1 (.I(_1550_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7338__I (.I(_2476_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7339__A1 (.I(_2467_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7339__B2 (.I(_2477_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7340__A1 (.I(_1678_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7340__A2 (.I(_1676_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7340__A3 (.I(_4240_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7341__I (.I(_2479_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7342__I (.I(_0853_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7343__I (.I(_2481_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7344__A1 (.I(_1463_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7344__A2 (.I(_2482_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7345__I (.I(_0885_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7346__A1 (.I(_2484_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7346__A2 (.I(_1311_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7347__I (.I(_2485_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7348__A1 (.I(_0863_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7348__A2 (.I(_4391_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7349__A1 (.I(_2486_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7349__A2 (.I(_2487_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7350__A1 (.I(_2418_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7350__A2 (.I(_2480_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7350__B (.I(_2483_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7351__A1 (.I(_1311_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7351__A2 (.I(_2478_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7352__A1 (.I(_1482_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7352__A2 (.I(_2481_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7353__I (.I(_2491_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7354__A1 (.I(_2150_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7354__A2 (.I(_4393_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7355__I (.I(_2493_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7356__I (.I(_2494_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7357__A1 (.I(_2492_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7357__A2 (.I(_2495_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7358__A2 (.I(_2487_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7359__A1 (.I(_2418_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7359__A2 (.I(_1710_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7360__A1 (.I(_0872_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7361__I (.I(_2499_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7362__A1 (.I(_2396_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7362__A2 (.I(_1684_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7364__I (.I(_0882_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7365__A1 (.I(_2153_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7365__A2 (.I(_2503_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7366__I (.I(_2504_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7367__A1 (.I(_0881_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7367__A2 (.I(_2154_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7368__I (.I(_2506_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7369__I (.I(_2507_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7370__I (.I(_2410_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7371__A1 (.I(_2417_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7371__A2 (.I(_2509_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7372__A1 (.I(_2418_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7372__A2 (.I(_2505_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7372__B1 (.I(_2508_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7372__B2 (.I(_1551_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7373__A2 (.I(_2500_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7373__B1 (.I(_2502_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7374__I (.I(_2492_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7375__I (.I(_1374_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7376__A1 (.I(_2145_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7376__A2 (.I(_2496_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7376__B1 (.I(_2512_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7376__B2 (.I(_2513_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7376__C (.I(_2514_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7377__A1 (.I(_2490_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7377__A2 (.I(_2515_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7377__B (.I(_2403_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7378__I (.I(_1359_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7379__A1 (.I(_0865_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7379__A2 (.I(_2517_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7379__B (.I(_2465_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7380__A1 (.I(_2418_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7380__A2 (.I(_2466_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7380__B1 (.I(_2516_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7381__A1 (.I(_2416_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7382__I (.I(_2464_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7383__I (.I(_2520_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7384__I (.I(_2517_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7385__A1 (.I(_1498_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7385__A2 (.I(_4418_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7386__I (.I(_2523_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7387__I (.I(_2524_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7388__A2 (.I(_2395_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7389__I (.I(_2526_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7390__A1 (.I(_2525_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7390__A2 (.I(_2527_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7391__A1 (.I(_1260_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7391__A2 (.I(_0872_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7393__A1 (.I(_2153_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7394__I (.I(_2531_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7395__I (.I(_0896_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7396__A1 (.I(_1340_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7396__A2 (.I(_2533_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7397__I (.I(_2534_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7398__I (.I(_4531_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7399__A1 (.I(_2530_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7399__A2 (.I(_2417_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7400__I (.I(_2154_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7401__I (.I(_2538_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7402__I (.I(_2539_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7403__A1 (.I(_2530_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7403__A2 (.I(_2532_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7403__B1 (.I(_2535_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7403__B2 (.I(_2536_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7403__C1 (.I(_2537_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7403__C2 (.I(_2540_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7404__I (.I(_1336_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7405__A1 (.I(\as2650.pc[0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7405__A2 (.I(net6));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7406__A1 (.I(_0910_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7406__A2 (.I(_4528_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7408__A1 (.I(_2542_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7408__A2 (.I(_2545_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7409__A1 (.I(_2530_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7409__A2 (.I(_1619_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7409__B (.I(_2499_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7410__A1 (.I(_2529_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7411__I (.I(_2523_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7412__I (.I(_2549_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7413__I (.I(_1569_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7414__A1 (.I(_0911_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7414__B2 (.I(_2550_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7414__C (.I(_2551_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7415__I (.I(_2469_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7416__I (.I(_1308_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7418__A1 (.I(_4390_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7418__A2 (.I(_4352_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7419__A1 (.I(_4529_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7419__A2 (.I(_0292_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7421__A1 (.I(_2536_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7421__A2 (.I(_2553_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7421__B (.I(_2554_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7422__I (.I(_2472_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7423__A1 (.I(_4390_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7424__A1 (.I(_4529_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7424__A2 (.I(_4513_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7427__I (.I(_2564_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7428__A1 (.I(_2536_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7428__C (.I(_2565_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7430__A1 (.I(_0862_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7430__A2 (.I(_4390_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7431__A1 (.I(_2568_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7432__I (.I(_1344_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7433__A1 (.I(_2486_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7433__A2 (.I(_2569_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7433__B (.I(_2570_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7434__A1 (.I(_2480_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7434__A2 (.I(_2537_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7434__B1 (.I(_2567_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7434__B2 (.I(_1337_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7435__I (.I(_1357_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7436__A2 (.I(_2572_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7437__A1 (.I(_0912_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7437__A2 (.I(_2522_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7438__A1 (.I(_2530_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7438__A2 (.I(_2520_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7439__I (.I(_1390_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7440__I (.I(_2577_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7441__A1 (.I(_2521_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7441__C (.I(_2578_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7442__I (.I(_2520_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7443__I (.I(_2517_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7444__I (.I(net7));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7445__A1 (.I(_0289_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7445__A2 (.I(_0291_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7445__B (.I(_2581_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7446__A1 (.I(_2581_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7446__A2 (.I(_0289_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7446__A3 (.I(_0291_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7448__B (.I(_0374_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7449__A1 (.I(_1554_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7449__A2 (.I(_0358_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7450__A1 (.I(_2585_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7451__I (.I(_4246_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7452__A1 (.I(_2584_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7452__B (.I(_2588_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7453__A1 (.I(_2584_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7454__A1 (.I(_1699_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7454__A2 (.I(_2553_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7454__B (.I(_2467_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7455__A1 (.I(_4503_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7455__A2 (.I(_0350_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7455__B1 (.I(_0356_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7455__B2 (.I(_0386_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7456__A1 (.I(_4511_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7456__A2 (.I(_4512_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7456__B (.I(_4528_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7457__A1 (.I(_4528_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7457__A2 (.I(_4511_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7457__A3 (.I(_4512_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7459__A1 (.I(_1553_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7459__A2 (.I(_2592_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7461__I (.I(_2564_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7462__A1 (.I(_1555_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7462__C (.I(_2598_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7464__A1 (.I(\as2650.pc[2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7464__A2 (.I(net8));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7466__A2 (.I(net7));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7467__A1 (.I(_0909_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7467__A2 (.I(net7));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7468__A1 (.I(_2568_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7470__I (.I(_1338_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7471__B (.I(_2607_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7473__A2 (.I(_2417_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7474__A1 (.I(_2609_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7475__I (.I(_1306_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7476__I (.I(_2612_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7477__A1 (.I(_2606_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7477__B1 (.I(_2611_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7477__B2 (.I(_2613_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7477__C (.I(_2570_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7478__A1 (.I(_1337_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7478__A2 (.I(_2600_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7479__A1 (.I(_2540_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7479__A2 (.I(_2611_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7480__A1 (.I(_2609_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7480__A2 (.I(_2505_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7480__B1 (.I(_2508_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7480__B2 (.I(_1555_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7481__I (.I(_2542_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7484__A2 (.I(_2620_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7485__A1 (.I(_2609_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7485__A2 (.I(_2618_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7485__B (.I(_2500_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7486__A1 (.I(_2529_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7487__I (.I(_1569_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7488__A1 (.I(_0921_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7488__B2 (.I(_2550_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7488__C (.I(_2624_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7489__A1 (.I(_2615_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7490__A1 (.I(_2178_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7490__A2 (.I(_2580_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7491__A1 (.I(_2609_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7491__A2 (.I(_2466_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7491__B (.I(_1635_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7492__A1 (.I(_2579_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7493__I (.I(_1283_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7494__I (.I(_2629_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7495__I (.I(_2443_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7496__I (.I(_2631_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7497__I (.I(_2632_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7498__I (.I(_1532_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7499__I (.I(_2634_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7500__A1 (.I(_2181_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7500__A2 (.I(_0506_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7501__A1 (.I(_0926_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7501__A2 (.I(_1584_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7502__A1 (.I(_2636_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7503__A1 (.I(\as2650.pc[2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7503__A2 (.I(_0373_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7505__A1 (.I(_2638_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7506__A1 (.I(_1614_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7506__A2 (.I(_2641_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7507__I (.I(net31));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7508__I (.I(_1579_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7509__I (.I(_2352_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7510__A1 (.I(_1684_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7510__A2 (.I(_2645_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7511__A1 (.I(_2643_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7511__A2 (.I(_2644_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7511__B (.I(_2646_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7514__A1 (.I(_2643_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7515__A1 (.I(_0508_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7515__A2 (.I(_1489_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7516__A1 (.I(_2648_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7516__A2 (.I(_2650_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7516__B1 (.I(_2651_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7516__B2 (.I(_1340_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7517__A1 (.I(_2643_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7517__A2 (.I(_2532_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7517__B (.I(_2652_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7518__B2 (.I(_2502_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7519__A1 (.I(_2335_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7519__A2 (.I(_2527_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7520__A1 (.I(_0928_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7520__A2 (.I(_2655_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7521__A1 (.I(_2635_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7521__A2 (.I(_2654_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7522__I (.I(_2340_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7523__A2 (.I(_2606_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7524__A1 (.I(_2638_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7525__A1 (.I(_2336_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7525__A2 (.I(_2479_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7526__I (.I(_1308_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7527__A1 (.I(_1585_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7527__A2 (.I(_0485_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7528__A1 (.I(_1584_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7530__A1 (.I(_0374_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7531__A1 (.I(_2584_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7531__A2 (.I(_2585_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7533__A1 (.I(_2469_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7533__A2 (.I(_2668_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7534__A1 (.I(_1594_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7534__B (.I(_2662_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7535__A1 (.I(_0375_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7535__A2 (.I(_2592_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7536__A1 (.I(_0374_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7536__A2 (.I(_2592_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7537__A2 (.I(_2672_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7538__A1 (.I(_1585_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7538__A2 (.I(_0491_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7539__A1 (.I(_2472_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7539__A2 (.I(_2674_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7540__A1 (.I(_1594_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7540__C (.I(_2564_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7542__A1 (.I(_2661_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7542__A2 (.I(_2677_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7542__B1 (.I(_2650_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7542__B2 (.I(_2479_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7542__C (.I(_2340_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7543__A1 (.I(_2658_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7543__A2 (.I(_2660_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7543__C (.I(_2483_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7544__A1 (.I(_0928_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7544__A2 (.I(_2630_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7544__B1 (.I(_2633_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7545__I (.I(_2403_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7546__A1 (.I(_2183_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7546__A2 (.I(_2580_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7546__B1 (.I(_2680_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7546__B2 (.I(_2681_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7547__A1 (.I(_2643_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7547__A2 (.I(_2466_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7547__B (.I(_1635_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7548__A1 (.I(_2579_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7549__I (.I(_2517_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7550__A1 (.I(_2190_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7550__A2 (.I(_2655_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7551__I (.I(_1513_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7553__I (.I(_2507_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7554__I (.I(net31));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7556__A1 (.I(_2687_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7556__A2 (.I(_2690_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7557__A1 (.I(_1582_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7557__A2 (.I(_2688_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7557__B1 (.I(_2691_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7557__B2 (.I(_2648_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7558__A1 (.I(_2687_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7558__A2 (.I(_2532_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7558__B (.I(_2502_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7559__I (.I(_0594_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7560__A1 (.I(_2187_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7560__A2 (.I(_2694_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7562__A1 (.I(_2636_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7563__A2 (.I(_2697_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7564__A2 (.I(_2698_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7565__A1 (.I(_2687_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7565__A2 (.I(_1710_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7565__B (.I(_2500_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7566__B (.I(_1252_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7567__A1 (.I(_2190_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7567__A2 (.I(_2686_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7567__B1 (.I(_1701_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7568__A1 (.I(\as2650.addr_buff[7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7569__I (.I(_2703_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7570__A1 (.I(_2565_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7570__A2 (.I(_2704_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7571__A1 (.I(_0507_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7571__A2 (.I(_0490_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7572__A1 (.I(_0507_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7572__A2 (.I(_0490_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7572__B2 (.I(_2672_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7573__A2 (.I(_2707_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7574__A1 (.I(_1581_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7574__A2 (.I(_0578_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7575__A1 (.I(_2584_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7575__A2 (.I(_2585_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7577__A2 (.I(_0614_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7578__A2 (.I(_2712_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7579__A1 (.I(_0597_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7579__A2 (.I(_2553_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7579__B (.I(_2554_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7580__A1 (.I(_1582_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7580__B1 (.I(_2709_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7580__B2 (.I(_4268_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7581__A1 (.I(_2181_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7581__A2 (.I(_0507_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7582__A1 (.I(_2636_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7584__I (.I(_2340_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7585__I (.I(_2612_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7586__A1 (.I(_2720_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7586__A2 (.I(_2691_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7586__B (.I(_2570_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7587__A1 (.I(_1337_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7587__A2 (.I(_2715_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7587__B1 (.I(_2718_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7587__B2 (.I(_2719_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7587__C (.I(_2721_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7588__B (.I(_2722_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7589__A1 (.I(_2191_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7589__A2 (.I(_2684_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7589__B1 (.I(_2723_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7589__B2 (.I(_2681_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7590__A1 (.I(_2687_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7590__A2 (.I(_2466_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7590__B (.I(_1635_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7591__A1 (.I(_2579_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7592__A1 (.I(_0939_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7592__A2 (.I(net1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7594__A1 (.I(_2188_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7594__A2 (.I(_0596_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7596__A1 (.I(_2728_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7596__A2 (.I(_2729_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7597__A1 (.I(_2727_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7598__A1 (.I(_0594_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7598__A2 (.I(_0613_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7599__A1 (.I(_2694_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7599__A2 (.I(_0613_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7601__A1 (.I(_1180_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7601__A2 (.I(_0668_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7602__I (.I(_0684_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7603__A1 (.I(_2736_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7603__A2 (.I(_4246_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7604__A1 (.I(_2588_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7604__A2 (.I(_2735_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7604__B (.I(_2737_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7604__C (.I(_2662_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7605__A1 (.I(_0595_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7605__A2 (.I(_0577_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7606__A1 (.I(_0595_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7606__A2 (.I(_0577_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7607__A3 (.I(_2707_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7608__A1 (.I(_1180_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7608__A2 (.I(_0698_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7608__A3 (.I(_2741_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7609__A1 (.I(_0685_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7609__A2 (.I(_2703_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7611__A1 (.I(_2704_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7611__A2 (.I(_2742_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7611__C (.I(_2744_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7613__A2 (.I(_2690_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7614__A1 (.I(net33));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7616__A1 (.I(_2661_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7616__A2 (.I(_2746_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7616__B1 (.I(_2749_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7616__B2 (.I(_2480_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7616__C (.I(_2658_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7617__I (.I(_2483_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7618__A1 (.I(_2719_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7618__C (.I(_2751_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7619__I (.I(_1701_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7620__I (.I(_2154_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7621__I (.I(_2754_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7622__I (.I(_2755_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7623__I (.I(net33));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7624__A1 (.I(_2757_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7624__A2 (.I(_2504_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7624__B1 (.I(_2688_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7624__B2 (.I(_2736_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7624__C (.I(_2529_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7625__A1 (.I(_2756_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7625__A2 (.I(_2749_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7626__A1 (.I(_0933_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7626__A2 (.I(_0594_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7627__A2 (.I(_2697_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7627__B (.I(_2728_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7628__A1 (.I(_2727_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7629__A1 (.I(_1680_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7629__A2 (.I(_2762_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7630__A1 (.I(_2757_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7630__A2 (.I(_1614_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7631__A1 (.I(_2499_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7633__A1 (.I(_0940_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7633__A2 (.I(_2655_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7633__B1 (.I(_2766_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7633__B2 (.I(_1443_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7634__A1 (.I(_2196_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7634__A2 (.I(_2686_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7634__B1 (.I(_2753_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7635__A1 (.I(_2752_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7636__A1 (.I(_2197_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7636__A2 (.I(_2580_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7637__I (.I(_2465_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7638__I (.I(_1634_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7639__A1 (.I(_2757_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7640__A1 (.I(_2579_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7641__I (.I(_2520_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7642__A1 (.I(_0948_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7642__A2 (.I(_2655_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7643__I (.I(_2503_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7644__I (.I(_2776_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7645__I (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7646__A1 (.I(_2757_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7647__A1 (.I(_2778_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7648__A1 (.I(_2778_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7648__A2 (.I(_2531_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7648__B1 (.I(_2534_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7648__B2 (.I(_1526_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7649__A1 (.I(_2777_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7649__A2 (.I(_2780_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7649__B (.I(_2781_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7650__A1 (.I(\as2650.pc[6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7650__A2 (.I(net2));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7652__A1 (.I(_2636_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7653__A1 (.I(_2194_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7653__A2 (.I(_0682_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7654__A1 (.I(_2194_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7654__A2 (.I(net1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7654__B (.I(net10));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7654__C (.I(_2187_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7656__A1 (.I(_2785_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7656__A2 (.I(_2788_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7658__A1 (.I(_2778_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7658__A2 (.I(_2542_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7658__B (.I(_2499_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7659__A1 (.I(_1619_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7659__A2 (.I(_2790_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7660__I (.I(_1271_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7661__I (.I(_2793_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7662__B (.I(_2794_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7663__A1 (.I(_2632_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7664__A1 (.I(_0948_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7664__A2 (.I(_2686_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7665__A1 (.I(_1587_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7665__A2 (.I(_0748_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7666__A1 (.I(_0682_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7666__A2 (.I(_0667_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7667__I (.I(_0682_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7668__A1 (.I(_2800_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7668__A2 (.I(_0667_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7672__A1 (.I(_1559_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7672__A2 (.I(_2553_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7672__B (.I(_2467_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7672__C (.I(_2804_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7673__A1 (.I(_1587_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7673__A2 (.I(_0770_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7674__A1 (.I(_2800_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7674__A2 (.I(_0697_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7675__A1 (.I(_0683_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7675__A2 (.I(_0697_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7676__A2 (.I(_2741_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7677__A2 (.I(_2809_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7679__A1 (.I(_1559_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7679__C (.I(_2565_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7680__B (.I(_1311_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7682__A1 (.I(_2729_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7682__A2 (.I(_2727_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7684__A2 (.I(_2816_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7685__I (.I(_2485_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7686__A1 (.I(_2613_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7686__A2 (.I(_2780_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7686__B2 (.I(_2818_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7687__A1 (.I(_2751_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7687__A2 (.I(_2813_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7689__A1 (.I(_2201_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7689__A2 (.I(_2684_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7689__B2 (.I(_2681_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7690__A1 (.I(_2778_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7691__A1 (.I(_2774_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7693__I (.I(_0756_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7694__A1 (.I(_2825_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7694__A2 (.I(_0749_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7696__A1 (.I(_1617_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7696__A2 (.I(_0828_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7697__A1 (.I(_1680_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7697__A2 (.I(_2588_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7698__A1 (.I(_2588_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7698__A2 (.I(_2828_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7698__C (.I(_2554_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7699__A1 (.I(_0757_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7699__A2 (.I(_0771_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7700__A2 (.I(_2809_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7701__A1 (.I(_1599_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7701__A2 (.I(_0830_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7702__A1 (.I(_1680_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7702__A2 (.I(_2704_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7703__A1 (.I(_2704_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7703__C (.I(_2476_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7705__B (.I(_2836_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7706__I (.I(net54));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7707__A1 (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7707__A2 (.I(net33));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7709__A1 (.I(_2720_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7709__B (.I(_2818_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7710__A1 (.I(\as2650.pc[7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7710__A2 (.I(net2));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7711__A1 (.I(_0945_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7711__A2 (.I(net2));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7712__A2 (.I(_2816_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7714__A1 (.I(_2837_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7714__B2 (.I(_2818_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7718__A1 (.I(_2618_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7718__A2 (.I(_2849_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7719__A1 (.I(_2491_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7719__A2 (.I(_2646_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7720__A1 (.I(_1516_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7721__A1 (.I(net54));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7721__A2 (.I(_2644_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7721__B (.I(_2852_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7722__I (.I(_1479_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7723__A1 (.I(_1497_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7723__A2 (.I(_1683_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7724__I (.I(_2855_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7725__A1 (.I(_2648_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7726__A1 (.I(net54));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7726__A2 (.I(_2505_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7726__B1 (.I(_2688_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7726__B2 (.I(_2542_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7727__A1 (.I(_2854_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7727__A2 (.I(_2856_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7728__A1 (.I(_2204_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7728__A2 (.I(_2496_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7729__B2 (.I(_1450_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7730__A1 (.I(_2751_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7731__A1 (.I(_2824_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7732__A1 (.I(_2205_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7732__A2 (.I(_2580_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7733__A1 (.I(net54));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7734__A1 (.I(_2774_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7736__A2 (.I(_0827_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7737__A1 (.I(_0836_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7737__A2 (.I(_0827_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7737__B (.I(_4245_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7738__I (.I(_2868_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7739__A1 (.I(_2866_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7739__A2 (.I(_2867_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7739__A3 (.I(_2869_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7740__I (.I(_2867_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7741__A1 (.I(_2871_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7741__A2 (.I(_2869_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7742__A1 (.I(_2334_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7744__A2 (.I(_0829_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7745__A2 (.I(_2809_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7746__A1 (.I(_1604_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7746__A2 (.I(_0829_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7747__A1 (.I(_2703_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7748__A1 (.I(_2866_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7748__A2 (.I(_2876_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7748__A3 (.I(_2878_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7749__A1 (.I(_2876_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7749__A2 (.I(_2878_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7750__A1 (.I(_2334_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7752__A1 (.I(_2467_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7752__A2 (.I(_2874_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7752__B1 (.I(_2882_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7752__B2 (.I(_2598_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7753__I (.I(net36));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7755__A1 (.I(_2884_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7755__A2 (.I(_2885_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7756__A1 (.I(_2480_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7756__A2 (.I(_2886_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7757__I (.I(_2485_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7758__A1 (.I(_2836_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7758__A2 (.I(_2883_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7758__C (.I(_2888_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7759__A1 (.I(\as2650.pc[8] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7761__A1 (.I(_2788_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7762__A1 (.I(_2203_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7763__A1 (.I(_2729_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7763__A2 (.I(_2727_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7765__B (.I(_2607_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7767__A1 (.I(_2895_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7767__B (.I(_2751_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7768__I (.I(_2866_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7769__A1 (.I(_2884_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7769__A2 (.I(_2532_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7769__B1 (.I(_2535_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7769__B2 (.I(_2899_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7769__C (.I(_2502_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7770__A1 (.I(_2386_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7770__A2 (.I(_2886_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7771__A1 (.I(_2785_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7773__A1 (.I(_2884_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7773__A2 (.I(_2618_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7773__B (.I(_2500_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7774__A1 (.I(_1546_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7774__A2 (.I(_2903_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7775__A1 (.I(_2901_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7775__B (.I(_2550_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7776__A1 (.I(_0966_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7776__B (.I(_2624_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7777__A1 (.I(_2889_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7778__A1 (.I(_0966_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7778__A2 (.I(_2684_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7778__B2 (.I(_2681_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7779__A1 (.I(_2884_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7780__A1 (.I(_2774_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7782__A2 (.I(_1586_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7783__A2 (.I(_0757_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7784__A2 (.I(_2895_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7786__A1 (.I(_2361_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7787__A1 (.I(_2361_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7788__A1 (.I(_2476_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7788__B2 (.I(_2554_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7789__I (.I(net37));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7790__A1 (.I(net36));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7790__A2 (.I(_2885_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7791__A1 (.I(_2919_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7792__A1 (.I(_2836_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7792__A2 (.I(_2918_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7792__B1 (.I(_2921_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7792__B2 (.I(_2720_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7792__C (.I(_2486_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7793__I (.I(_2570_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7794__A1 (.I(_2818_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7794__B (.I(_2922_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7794__C (.I(_2923_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7795__I (.I(_1479_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7796__I (.I(_2925_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7797__I (.I(_2855_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7798__I (.I(_2927_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7799__A1 (.I(_2777_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7799__A2 (.I(_2921_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7800__A1 (.I(_2919_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7800__A2 (.I(_2505_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7800__B1 (.I(_2688_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7800__B2 (.I(_2362_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7801__A1 (.I(_2926_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7801__A2 (.I(_2928_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7802__A1 (.I(_0979_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7802__A2 (.I(_2496_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7803__A1 (.I(_2514_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7807__A1 (.I(_2919_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7807__A2 (.I(_2644_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7807__B (.I(_2852_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7808__A1 (.I(_2377_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7810__I (.I(_1327_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7811__A1 (.I(_0979_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7811__A2 (.I(_2684_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7811__B2 (.I(_2940_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7812__I (.I(_2465_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7813__I (.I(_1565_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7814__A1 (.I(_2919_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7814__A2 (.I(_2942_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7814__B (.I(_2943_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7815__A1 (.I(_2774_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7816__I (.I(net53));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7817__A1 (.I(net37));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7817__A2 (.I(net36));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7817__A3 (.I(_2885_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7819__A1 (.I(_2744_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7819__A2 (.I(_2876_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7819__A3 (.I(_2878_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7820__A1 (.I(_2662_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7820__A2 (.I(_2871_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7820__A3 (.I(_2869_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7821__A1 (.I(_2899_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7821__A2 (.I(_2361_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7821__A3 (.I(_2366_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7822__B (.I(_2950_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7823__A1 (.I(_2866_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7823__A2 (.I(\as2650.addr_buff[1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7824__A1 (.I(_2871_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7824__A2 (.I(_2869_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7824__B (.I(_2564_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7825__A1 (.I(_2336_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7825__A2 (.I(_2612_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7825__B1 (.I(_2952_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7826__A2 (.I(_2952_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7826__B (.I(_2744_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7827__B (.I(_2366_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7828__B (.I(_2661_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7829__A1 (.I(_2613_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7829__B (.I(_2957_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7829__C (.I(_2888_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7830__A2 (.I(_1586_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7832__B (.I(_0756_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7833__I (.I(_2961_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7834__A1 (.I(_2895_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7835__A3 (.I(_2963_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7836__A2 (.I(_2963_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7837__A1 (.I(_2658_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7838__A1 (.I(_2923_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7841__A1 (.I(_2540_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7842__A1 (.I(net53));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7842__A2 (.I(_2531_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7842__B1 (.I(_2535_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7842__B2 (.I(_2366_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7842__C (.I(_2854_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7843__A1 (.I(_2969_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7843__A2 (.I(_2527_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7843__B2 (.I(_2971_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7844__A1 (.I(_0990_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7844__A2 (.I(_2513_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7844__B2 (.I(_2928_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7844__C (.I(_2551_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7846__A1 (.I(_2961_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7846__A2 (.I(_2974_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7848__A1 (.I(_1546_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7848__A2 (.I(_2976_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7849__A1 (.I(net53));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7849__A2 (.I(_1711_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7850__A2 (.I(_2967_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7851__A1 (.I(_0990_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7851__A2 (.I(_2522_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7851__B2 (.I(_2940_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7852__A1 (.I(net53));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7852__A2 (.I(_2942_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7852__B (.I(_2943_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7853__A1 (.I(_2521_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7854__I (.I(net39));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7856__A1 (.I(_2982_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7857__A2 (.I(_2950_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7857__B (.I(_2612_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7858__A2 (.I(_2950_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7858__B (.I(_2744_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7859__A1 (.I(_2369_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7860__A1 (.I(_2369_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7860__C (.I(_2661_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7861__A1 (.I(_2613_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7861__A2 (.I(_2984_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7861__B (.I(_2988_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7861__C (.I(_2888_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7862__A1 (.I(\as2650.pc[11] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7862__A2 (.I(_1586_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7863__A1 (.I(_0989_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7863__A2 (.I(_0757_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7866__A1 (.I(_2719_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7866__A2 (.I(_2993_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7866__B (.I(_2483_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7867__I (.I(_0997_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7868__I (.I(_2494_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7869__A1 (.I(_2385_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7869__A2 (.I(_2984_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7870__I (.I(\as2650.addr_buff[3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7871__A1 (.I(_2982_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7871__A2 (.I(_2504_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7871__B1 (.I(_2507_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7871__B2 (.I(_2998_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7871__C (.I(_1268_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7872__A1 (.I(_2995_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7872__A2 (.I(_2996_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7873__I (.I(_2149_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7874__A1 (.I(_0997_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7874__A2 (.I(_2525_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7874__B2 (.I(_3001_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7875__A1 (.I(_1575_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7879__A1 (.I(_2982_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7879__A2 (.I(_2644_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7880__A1 (.I(_1546_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7880__A2 (.I(_3006_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7880__C (.I(_2852_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7882__A1 (.I(_0997_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7882__A2 (.I(_2522_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7882__B2 (.I(_2940_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7883__A1 (.I(_2982_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7883__A2 (.I(_2942_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7883__B (.I(_2943_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7884__A1 (.I(_2521_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7885__A1 (.I(\as2650.pc[12] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7885__A2 (.I(_0756_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7888__A1 (.I(\as2650.pc[11] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7888__B (.I(_2825_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7889__A1 (.I(_2974_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7889__C (.I(_2961_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7891__A1 (.I(_1711_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7891__A2 (.I(_3017_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7892__A1 (.I(net52));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7892__A2 (.I(_2377_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7892__B (.I(_2852_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7893__I (.I(\as2650.addr_buff[4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7894__A2 (.I(\as2650.addr_buff[1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7895__A1 (.I(_2998_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7895__A2 (.I(_2871_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7895__A3 (.I(_2868_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7895__A4 (.I(_3021_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7896__A1 (.I(_3020_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7897__A1 (.I(_2998_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7897__A2 (.I(_2876_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7897__A3 (.I(_2878_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7897__A4 (.I(_3021_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7898__A1 (.I(_3020_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7899__A1 (.I(_2662_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7899__B2 (.I(_2476_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7900__A1 (.I(net39));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7901__A1 (.I(net52));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7902__A1 (.I(_2836_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7902__A2 (.I(_3026_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7902__B1 (.I(_3028_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7902__B2 (.I(_2720_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7902__C (.I(_2486_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7903__A1 (.I(_2961_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7904__A1 (.I(_2963_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7906__A1 (.I(_2607_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7906__A2 (.I(_3032_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7907__A1 (.I(_2923_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7907__A2 (.I(_3029_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7908__I (.I(\as2650.pc[12] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7909__A1 (.I(_2385_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7909__A2 (.I(_3028_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7910__A1 (.I(net52));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7910__A2 (.I(_2504_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7910__B1 (.I(_2507_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7910__B2 (.I(_3020_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7910__C (.I(_1268_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7911__A1 (.I(_3035_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7911__A2 (.I(_2495_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7912__A1 (.I(_1003_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7912__A2 (.I(_2525_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7912__B2 (.I(_3001_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7913__A1 (.I(_1450_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7914__A1 (.I(_3018_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7915__A1 (.I(_1003_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7915__A2 (.I(_2522_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7915__B2 (.I(_2940_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7916__A1 (.I(net52));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7916__A2 (.I(_2942_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7916__B (.I(_2943_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7917__A1 (.I(_2521_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7918__I (.I(_2445_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7919__I (.I(_1320_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7920__A1 (.I(_1462_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7920__A2 (.I(_1327_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7921__A1 (.I(_3045_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7921__A2 (.I(_2354_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7921__A3 (.I(_3046_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7921__A4 (.I(_2433_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7922__I (.I(_0871_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7923__A1 (.I(_3048_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7923__A2 (.I(_2152_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7923__B (.I(_4444_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7924__A1 (.I(_1331_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7924__A2 (.I(_2412_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7925__A1 (.I(_1480_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7925__A2 (.I(_2427_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7926__A2 (.I(_2425_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7927__A1 (.I(_4491_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7927__A2 (.I(_2446_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7928__A1 (.I(_1353_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7928__A2 (.I(_3050_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7928__A3 (.I(_3052_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7928__A4 (.I(_3053_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7929__A1 (.I(_2422_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7929__A2 (.I(_2453_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7930__A4 (.I(_3055_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7931__I (.I(_2157_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7933__I (.I(_3058_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7934__A1 (.I(_2551_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7934__A2 (.I(_4187_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7934__A3 (.I(_3059_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7935__I (.I(_1324_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7936__A1 (.I(net26));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7936__A2 (.I(_1367_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7936__B1 (.I(_3061_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7936__B2 (.I(_1575_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7936__C (.I(_1443_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7937__A1 (.I(_2686_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7937__A2 (.I(_2381_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7937__B1 (.I(_3060_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7938__A1 (.I(_2824_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7938__A2 (.I(_3063_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7938__B (.I(_3056_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7939__A2 (.I(_3056_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7939__C (.I(_2578_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7940__A1 (.I(_1356_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7940__A2 (.I(_1684_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7940__A3 (.I(_1504_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7941__A2 (.I(_2348_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7942__A1 (.I(_0891_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7943__A1 (.I(_3065_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7943__A2 (.I(_3067_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7944__A1 (.I(_2349_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7946__A1 (.I(_4237_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7946__A2 (.I(_2348_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7946__A3 (.I(_3070_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7947__A1 (.I(_3069_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7947__A2 (.I(_3071_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7948__A1 (.I(_4490_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7948__A2 (.I(_2444_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7948__A3 (.I(_2446_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7949__I (.I(_1503_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7950__A1 (.I(_2450_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7950__A2 (.I(_3074_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7950__A3 (.I(_2412_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7950__A4 (.I(_2451_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7951__I (.I(_2157_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7952__A1 (.I(_2396_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7952__A2 (.I(_3076_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7952__B1 (.I(_2407_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7952__B2 (.I(_1163_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7952__C (.I(_1319_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7953__A1 (.I(_1087_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7953__A2 (.I(_2441_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7954__A2 (.I(_3075_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7955__I (.I(_1516_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7956__A1 (.I(_1617_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7956__A2 (.I(_2352_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7957__I (.I(_2493_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7958__A1 (.I(_1482_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7958__A2 (.I(_1293_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7958__A3 (.I(_2160_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7958__A4 (.I(_3082_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7959__A1 (.I(_2149_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7959__A2 (.I(_3081_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7960__A1 (.I(_3080_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7962__A1 (.I(_2463_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7963__I (.I(_1517_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7964__I (.I(_1275_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7965__I (.I(_3089_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7966__A1 (.I(net51));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7966__A2 (.I(_3090_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7967__A1 (.I(_2380_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7967__B (.I(_1481_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7968__I (.I(_2160_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7969__A1 (.I(_3093_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7969__A2 (.I(_2155_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7969__B (.I(_2508_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7970__I (.I(_0872_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7971__A1 (.I(net51));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7971__A2 (.I(_1277_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7971__A3 (.I(_3095_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7972__C (.I(_2525_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7973__A2 (.I(_3097_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7974__A1 (.I(net51));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7974__A2 (.I(_3090_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7974__A3 (.I(_2155_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7975__A1 (.I(_3088_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7975__B2 (.I(_2923_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7976__A1 (.I(_1692_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7976__B (.I(_2403_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7977__A1 (.I(net51));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7977__A2 (.I(_3087_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7978__A1 (.I(_3087_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7978__C (.I(_2578_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7979__I (.I(_2793_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7980__A1 (.I(_3103_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7980__A2 (.I(_2338_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7980__A3 (.I(_1312_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7981__A1 (.I(_2551_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7982__I (.I(_1486_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7983__A1 (.I(_2407_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7983__C (.I(_3106_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7984__A1 (.I(_4265_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7984__A2 (.I(_2824_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7985__A2 (.I(_3107_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7986__A1 (.I(_3107_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7986__C (.I(_2578_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7987__A1 (.I(_4264_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7987__A2 (.I(_2824_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7988__A2 (.I(_3107_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7989__I (.I(_2577_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7990__A1 (.I(_3107_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7990__C (.I(_3112_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7991__A1 (.I(_4406_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7991__A2 (.I(_1524_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7992__A1 (.I(_1550_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7992__A2 (.I(_1442_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7993__A1 (.I(_3113_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7993__A2 (.I(_3114_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7994__A1 (.I(_1367_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7994__A2 (.I(_2420_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7995__A1 (.I(_1457_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7995__A2 (.I(_1477_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7995__B (.I(_1571_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7996__A1 (.I(_1277_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7996__A2 (.I(_1493_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7996__B (.I(_1517_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7996__C (.I(_0852_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7998__I (.I(_3119_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7999__I0 (.I(_3115_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7999__I1 (.I(_4291_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7999__S (.I(_3120_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8001__A1 (.I(_2536_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8001__A2 (.I(_1289_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8002__A1 (.I(_4542_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8002__A2 (.I(_1294_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8003__A1 (.I(_3122_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8003__A2 (.I(_3123_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8004__I0 (.I(_3124_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8004__I1 (.I(_0297_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8004__S (.I(_3120_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8006__I (.I(_1289_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8007__A1 (.I(_0361_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8007__A2 (.I(_3126_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8008__A1 (.I(_1699_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8008__A2 (.I(_1295_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8010__I (.I(_3119_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8011__I0 (.I(_3129_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8011__I1 (.I(_0413_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8011__S (.I(_3130_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8013__A1 (.I(_1594_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8013__A2 (.I(_1622_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8014__A1 (.I(_0535_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8014__A2 (.I(_1295_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8014__B (.I(_3132_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8015__A1 (.I(_0461_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8015__A2 (.I(_3120_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8016__A1 (.I(_3120_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8016__A2 (.I(_3133_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8017__A1 (.I(_0579_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8017__A2 (.I(_2399_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8018__I (.I(_2794_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8019__A1 (.I(_1558_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8019__A2 (.I(_3136_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8021__I0 (.I(_3138_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8021__I1 (.I(_0549_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8021__S (.I(_3130_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8023__A1 (.I(_2736_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8023__A2 (.I(_3103_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8024__A1 (.I(_1290_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8024__A2 (.I(_3140_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8025__I0 (.I(_3141_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8025__I1 (.I(_0637_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8025__S (.I(_3130_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8027__I (.I(_1524_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8028__I (.I(_3143_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8029__A1 (.I(_1706_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8029__A2 (.I(_1572_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8030__A1 (.I(_1530_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8030__A2 (.I(_3144_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8031__I0 (.I(_3146_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8031__S (.I(_3130_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8033__A1 (.I(_1710_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8033__A2 (.I(_1294_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8034__A2 (.I(_3148_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8035__I0 (.I(_3149_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8035__S (.I(_3119_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8037__A1 (.I(_2416_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8037__A2 (.I(_1488_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8038__I (.I(_3106_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8039__A1 (.I(_3151_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8039__A2 (.I(_1677_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8040__I (.I(_1685_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8041__I (.I(_2149_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8042__A1 (.I(_2440_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8042__A2 (.I(_2461_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8043__A1 (.I(_1250_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8043__A2 (.I(_3155_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8044__I (.I(_2503_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8045__I (.I(_3157_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8046__A1 (.I(_1676_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8046__A2 (.I(_1268_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8047__A1 (.I(_3158_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8048__A1 (.I(_3156_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8048__B (.I(_3059_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8049__A1 (.I(_1354_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8049__A2 (.I(_2348_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8050__I (.I(_0898_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8051__I (.I(_3163_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8052__A1 (.I(_2535_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8052__A2 (.I(_3162_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8052__B (.I(_3164_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8053__A1 (.I(_1237_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8053__A2 (.I(_1045_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8053__A3 (.I(_1273_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8054__A1 (.I(_1676_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8054__A2 (.I(_1236_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8054__A3 (.I(_1249_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8055__A1 (.I(_3158_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8055__A2 (.I(_1370_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8055__B2 (.I(_3167_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8056__A1 (.I(_1612_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8056__A2 (.I(_1256_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8056__B (.I(_1229_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8056__C (.I(_2482_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8057__I (.I(_3045_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8058__A1 (.I(_1249_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8058__B (.I(_3169_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8058__C (.I(_3170_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8060__A1 (.I(_3154_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8060__A3 (.I(_3165_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8060__B (.I(_3172_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8061__A1 (.I(_1677_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8061__A2 (.I(_3153_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8061__B1 (.I(_2407_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8062__I (.I(_4241_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8063__A1 (.I(_2618_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8063__A2 (.I(_0687_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8063__B (.I(_2607_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8064__A1 (.I(_1354_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8064__A2 (.I(_3175_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8064__B (.I(_2390_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8065__I (.I(_1342_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8066__A1 (.I(_0687_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8066__A2 (.I(_3175_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8067__A1 (.I(_3178_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8069__A1 (.I(_1272_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8069__A2 (.I(_3181_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8071__I (.I(_3183_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8072__A3 (.I(_3184_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8073__A1 (.I(_4417_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8073__A2 (.I(_1279_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8074__A2 (.I(_3186_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8075__A1 (.I(_1570_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8075__A2 (.I(_3174_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8075__B1 (.I(_3185_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8075__B2 (.I(_3187_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8075__C (.I(_2400_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8076__I (.I(_1391_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8077__B (.I(_3189_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8078__A1 (.I(_3151_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8078__A2 (.I(_1678_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8079__I (.I(_1498_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8081__A1 (.I(_3191_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8081__A2 (.I(_3192_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8081__B1 (.I(_3067_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8081__B2 (.I(_3154_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8082__I (.I(_1685_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8083__A1 (.I(_2383_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8083__A2 (.I(_3061_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8083__A3 (.I(_3192_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8084__A1 (.I(_3194_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8084__A2 (.I(_3156_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8084__B (.I(_3195_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8085__A1 (.I(_3164_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8086__A1 (.I(_2399_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8086__A2 (.I(_3167_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8087__I (.I(_3170_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8088__A1 (.I(_2383_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8088__A2 (.I(_3192_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8088__B (.I(_3169_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8088__C (.I(_3199_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8089__C (.I(_2624_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8090__A1 (.I(_3178_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8090__A2 (.I(_3192_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8091__A1 (.I(_2888_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8092__A1 (.I(_3136_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8092__A2 (.I(_3061_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8093__A1 (.I(_3186_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8093__A2 (.I(_3204_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8093__B (.I(_1576_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8094__A1 (.I(_3201_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8094__B (.I(_4201_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8095__B (.I(_3189_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8096__I (.I(_3106_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8097__I (.I(_3207_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8099__I (.I(_3046_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8100__A1 (.I(_2386_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8100__A2 (.I(_3090_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8100__B (.I(_1370_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8101__A1 (.I(_3209_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8101__A2 (.I(_1507_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8102__A1 (.I(_3090_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8102__A2 (.I(_1231_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8102__B (.I(_3212_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8103__I (.I(_3045_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8104__A1 (.I(_1304_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8104__A2 (.I(_4175_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8104__B (.I(_3214_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8105__I (.I(_2388_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8106__A1 (.I(_3211_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8107__A1 (.I(_3211_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8107__B2 (.I(_3216_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8108__I (.I(_3158_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8109__A1 (.I(_3219_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8109__A2 (.I(_3212_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8111__A1 (.I(_3164_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8111__A2 (.I(_3221_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8111__B (.I(_3067_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8112__A1 (.I(_4253_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8112__A2 (.I(_3153_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8112__B1 (.I(_2508_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8112__B2 (.I(_3059_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8112__C (.I(_3191_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8113__A1 (.I(_3220_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8113__A2 (.I(_3222_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8114__A1 (.I(_3210_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8115__I (.I(_1328_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8116__A1 (.I(_1429_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8116__A2 (.I(_1493_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8116__B (.I(_3220_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8117__A1 (.I(_3226_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8117__A2 (.I(_3227_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8117__B (.I(_3207_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8118__I (.I(_1301_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8119__A1 (.I(_3208_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8119__A2 (.I(_3209_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8119__B1 (.I(_3225_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8119__C (.I(_3229_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8120__I (.I(_3170_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8121__A1 (.I(_1681_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8121__A2 (.I(_2155_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8121__B (.I(_3221_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8122__A1 (.I(_3209_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8122__A2 (.I(_1507_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8123__A1 (.I(_0893_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8124__A1 (.I(_3230_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8124__A2 (.I(_3231_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8125__A1 (.I(_1451_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8126__A1 (.I(_0869_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8126__A2 (.I(_2506_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8127__A1 (.I(_3081_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8127__A2 (.I(_3236_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8129__A1 (.I(_0687_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8129__A2 (.I(_2658_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8129__B1 (.I(_3178_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8130__A1 (.I(_2624_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8130__A2 (.I(_3061_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8130__A3 (.I(_1339_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8130__A4 (.I(_2390_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8131__B (.I(_4201_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8132__A1 (.I(_2633_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8132__A2 (.I(_3237_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8133__A1 (.I(_3151_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8133__A2 (.I(_0893_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8133__C (.I(_3229_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8135__A1 (.I(_1486_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8135__A2 (.I(_0893_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8135__A3 (.I(_3209_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8135__A4 (.I(_1507_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8136__I (.I(_1565_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8137__B (.I(_3245_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8141__A1 (.I(_2416_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8142__I (.I(_1301_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8143__I (.I(_4171_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8144__A1 (.I(_2150_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8144__A2 (.I(_3250_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8144__B (.I(_1339_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8144__C (.I(_3178_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8145__A3 (.I(\as2650.cycle[3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8146__A1 (.I(_2484_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8146__A2 (.I(_3252_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8147__A1 (.I(_3175_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8147__A2 (.I(_3226_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8148__A1 (.I(_3226_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8148__A2 (.I(_3251_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8148__C (.I(_3207_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8149__A1 (.I(_3208_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8149__A2 (.I(_2484_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8149__B (.I(_3249_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8151__I (.I(_3256_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8152__A1 (.I(_1572_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8152__A2 (.I(_2477_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8152__A3 (.I(_2719_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8152__B (.I(_3226_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8153__A1 (.I(_2484_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8153__A2 (.I(_3252_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8154__A1 (.I(_1329_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8155__A1 (.I(_1570_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8155__A2 (.I(_3257_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8155__C (.I(_3207_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8156__A1 (.I(_3208_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8156__A2 (.I(_1329_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8156__B (.I(_3229_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8157__I (.I(\as2650.psu[7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8159__A1 (.I(_3263_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8159__A2 (.I(_3074_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8160__I (.I(_4420_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8161__A1 (.I(_3265_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8161__A2 (.I(_1527_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8162__A1 (.I(_1711_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8162__A2 (.I(_3266_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8163__A1 (.I(_4176_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8163__A2 (.I(_1510_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8164__A1 (.I(\as2650.psu[7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8164__A2 (.I(_2377_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8164__B (.I(_3268_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8165__A1 (.I(_0791_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8165__A2 (.I(_3074_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8167__A2 (.I(_3271_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8167__B (.I(_3151_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8168__A1 (.I(_3262_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8168__A2 (.I(_3208_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8168__B (.I(_3229_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8168__C (.I(_3272_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8169__A1 (.I(_0867_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8169__A2 (.I(_0879_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8169__A3 (.I(_1682_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8169__A4 (.I(_2346_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8170__A1 (.I(_3236_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8170__A2 (.I(_3273_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8171__A1 (.I(_2439_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8171__A2 (.I(_3186_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8172__A1 (.I(_0853_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8172__A2 (.I(_1248_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8172__A3 (.I(_2427_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8173__A1 (.I(_2428_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8174__A1 (.I(_2631_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8175__A1 (.I(_2336_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8175__A2 (.I(_0885_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8175__A3 (.I(_1462_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8176__A1 (.I(_2156_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8176__A2 (.I(_2506_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8176__B (.I(_1364_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8176__C (.I(_4200_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8177__A1 (.I(_1322_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8177__A2 (.I(_0889_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8177__C (.I(_3280_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8178__A1 (.I(_1347_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8178__A2 (.I(_1363_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8179__A1 (.I(_4444_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8179__A2 (.I(_2435_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8179__A3 (.I(_3281_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8180__A3 (.I(_3283_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8181__A1 (.I(_3157_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8181__A2 (.I(_3163_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8181__A3 (.I(_1349_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8181__A4 (.I(_3065_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8182__A1 (.I(_3052_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8182__A2 (.I(_3069_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8182__A3 (.I(_3071_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8183__A1 (.I(_3055_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8183__A3 (.I(_3285_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8184__I (.I(_3287_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8185__I (.I(_3288_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8186__I (.I(_1358_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8187__I (.I(_3290_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8188__I (.I(_3291_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8189__I (.I(_3095_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8190__A2 (.I(_1605_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8191__A1 (.I(_1544_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8191__A2 (.I(_2487_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8193__C (.I(_1509_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8194__A1 (.I(_4392_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8194__A2 (.I(_2410_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8195__A1 (.I(_2899_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8195__A2 (.I(_2755_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8195__B (.I(_1276_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8196__A1 (.I(_1442_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8196__A3 (.I(_3299_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8197__A1 (.I(\as2650.pc[0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8197__A2 (.I(_4180_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8198__A2 (.I(_3301_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8199__A1 (.I(_2458_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8199__A2 (.I(_0834_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8200__I0 (.I(_2145_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8200__S (.I(_3303_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8201__A1 (.I(_2440_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8202__A1 (.I(_0864_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8202__A2 (.I(_2440_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8202__C (.I(_4161_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8203__A1 (.I(_4161_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8203__C (.I(_1251_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8204__A1 (.I(_3093_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8205__A1 (.I(_2754_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8205__A2 (.I(_4281_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8206__A1 (.I(_1549_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8207__A1 (.I(_2382_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8207__A2 (.I(_3310_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8208__A1 (.I(_0864_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8208__A2 (.I(_2854_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8208__B (.I(_3058_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8209__A1 (.I(_3293_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8210__A1 (.I(_2335_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8211__A1 (.I(_2145_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8211__A2 (.I(_2794_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8211__B (.I(_3194_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8212__A1 (.I(_3214_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8213__I (.I(_2387_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8214__A1 (.I(\as2650.stack[7][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8214__A2 (.I(_1919_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8214__B1 (.I(_1638_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8215__I (.I(_1902_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8216__I (.I(_1654_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8217__A1 (.I(\as2650.stack[4][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8217__A2 (.I(_3319_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8217__B2 (.I(\as2650.stack[5][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8217__C (.I(_4475_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8218__I (.I(_1637_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8219__A1 (.I(\as2650.stack[3][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8219__A2 (.I(_1918_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8219__B1 (.I(_1902_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8219__C1 (.I(\as2650.stack[1][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8219__C2 (.I(_1654_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8221__A1 (.I(\as2650.stack[2][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8221__A2 (.I(_3322_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8221__B (.I(_0328_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8223__I (.I(_2408_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8224__A1 (.I(_0864_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8224__A2 (.I(_3317_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8224__B1 (.I(_3326_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8224__B2 (.I(_3327_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8225__I (.I(_3290_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8226__A1 (.I(_3316_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8226__B (.I(_3329_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8227__I (.I(_3287_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8228__A1 (.I(_0865_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8228__A2 (.I(_3292_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8228__C (.I(_3331_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8229__A1 (.I(_0865_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8229__A2 (.I(_3289_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8229__C (.I(_3112_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8230__I (.I(_3291_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8231__A1 (.I(_0910_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8233__I (.I(_2387_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8234__A1 (.I(_3336_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8234__A2 (.I(_3335_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8235__A1 (.I(_1677_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8235__A2 (.I(_3335_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8235__B (.I(_2926_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8236__A1 (.I(net6));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8236__A2 (.I(_4281_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8237__A1 (.I(_4530_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8237__A2 (.I(_4380_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8238__A1 (.I(_4530_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8238__A2 (.I(_2503_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8239__A1 (.I(_2777_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8239__C (.I(_3089_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8240__A1 (.I(_1696_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8240__A2 (.I(_1681_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8240__A3 (.I(_3342_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8241__A1 (.I(_2362_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8241__A2 (.I(_3181_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8242__I (.I(_2533_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8243__A1 (.I(_4531_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8243__A2 (.I(_3345_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8244__A1 (.I(_3089_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8244__A2 (.I(_2438_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8245__A1 (.I(_1696_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8245__B (.I(_1276_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8246__A1 (.I(_1679_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8246__A2 (.I(_2545_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8247__A1 (.I(_0911_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8247__A2 (.I(_1618_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8248__A1 (.I(_3048_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8248__B1 (.I(_3350_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8248__B2 (.I(_1696_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8249__A1 (.I(_2335_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8250__I (.I(_3155_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8251__A1 (.I(_1681_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8251__A2 (.I(_3353_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8252__A1 (.I(_0909_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8252__A2 (.I(_3301_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8253__A1 (.I(_0911_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8253__A2 (.I(_3301_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8254__A1 (.I(_3355_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8255__A2 (.I(_3335_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8255__C (.I(_1289_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8256__A2 (.I(_3343_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8257__A2 (.I(_4474_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8257__B (.I(_4473_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8260__A2 (.I(_1637_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8261__A2 (.I(_3361_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8261__B1 (.I(_3362_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8261__B2 (.I(\as2650.stack[1][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8262__A2 (.I(_3361_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8262__B1 (.I(_3362_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8262__B2 (.I(\as2650.stack[5][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8263__I (.I(_1918_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8264__A2 (.I(_3366_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8264__B1 (.I(_3322_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8264__C (.I(_4476_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8265__A1 (.I(_3360_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8266__I (.I(_2391_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8267__A1 (.I(_3199_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8267__B1 (.I(_3368_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8267__B2 (.I(_3369_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8268__I (.I(_3290_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8269__A2 (.I(_3370_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8269__B (.I(_3371_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8270__I (.I(_3287_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8271__I (.I(_3373_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8272__A1 (.I(_3333_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8272__A2 (.I(_3335_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8272__C (.I(_3374_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8273__A1 (.I(_3055_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8273__A3 (.I(_3285_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8274__I (.I(_3376_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8275__A1 (.I(_2170_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8275__A2 (.I(_3377_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8275__B (.I(_1566_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8277__I (.I(_3291_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8278__A1 (.I(_0910_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8278__A2 (.I(_0862_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8279__A1 (.I(_0919_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8281__A2 (.I(_4474_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8281__B (.I(_4473_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8282__A2 (.I(_3322_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8283__A2 (.I(_3319_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8283__B2 (.I(\as2650.stack[1][2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8284__I (.I(_1637_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8285__A2 (.I(_1918_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8285__B1 (.I(_1902_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8285__B2 (.I(\as2650.stack[4][2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8285__C1 (.I(\as2650.stack[5][2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8285__C2 (.I(_1654_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8286__A1 (.I(_0327_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8287__A2 (.I(_3386_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8288__A3 (.I(_3385_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8289__I (.I(_3095_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8290__A1 (.I(_1267_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8290__B1 (.I(_3155_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8290__B2 (.I(_1288_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8291__I (.I(_3392_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8292__A1 (.I(_1271_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8292__A2 (.I(_2157_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8292__A3 (.I(_3155_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8293__I (.I(_3394_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8294__A2 (.I(_3355_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8295__A1 (.I(_3395_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8296__A1 (.I(_3382_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8296__A2 (.I(_3393_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8296__B (.I(_3397_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8297__A1 (.I(_0373_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8297__A2 (.I(_4517_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8298__A1 (.I(_1553_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8298__A2 (.I(_4517_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8300__A1 (.I(_2581_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8300__A2 (.I(_4380_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8301__A1 (.I(_2581_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8301__A2 (.I(_4380_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8304__A1 (.I(_1553_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8304__A2 (.I(_2538_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8305__A1 (.I(_2509_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8305__B (.I(_3406_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8306__A1 (.I(_0919_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8306__A2 (.I(_1708_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8307__A1 (.I(_1336_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8307__A2 (.I(_2620_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8308__A1 (.I(_2365_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8308__A2 (.I(_2754_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8309__A1 (.I(_0376_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8309__A2 (.I(_2533_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8309__B (.I(_1508_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8310__A1 (.I(_3082_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8310__B1 (.I(_3409_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8310__B2 (.I(_2645_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8310__C (.I(_3411_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8311__A1 (.I(_3093_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8312__A1 (.I(_3070_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8312__A2 (.I(_3407_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8314__A1 (.I(_3415_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8314__A2 (.I(_3382_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8314__B1 (.I(_3409_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8314__B2 (.I(_2549_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8314__C (.I(_2856_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8315__A1 (.I(_3391_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8315__B1 (.I(_3414_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8315__B2 (.I(_2345_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8316__A1 (.I(_3336_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8316__A2 (.I(_3382_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8316__B1 (.I(_3390_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8316__B2 (.I(_3369_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8317__A1 (.I(_3329_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8317__A2 (.I(_3382_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8318__I (.I(_3376_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8319__A1 (.I(_3379_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8319__C (.I(_3420_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8320__A1 (.I(_2178_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8320__A2 (.I(_3377_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8321__A1 (.I(_2416_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8321__A2 (.I(_3422_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8322__A1 (.I(\as2650.pc[2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8322__A2 (.I(_0909_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8322__A3 (.I(\as2650.pc[0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8323__A2 (.I(_3423_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8324__I (.I(_3424_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8325__I (.I(_2387_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8326__A1 (.I(_2181_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8326__A2 (.I(_0919_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8326__A3 (.I(_3355_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8328__A2 (.I(_3355_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8328__B (.I(_2182_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8329__A1 (.I(_1293_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8329__A2 (.I(_3353_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8330__A1 (.I(_3428_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8330__A2 (.I(_3429_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8331__A1 (.I(_2182_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8331__A2 (.I(_1617_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8332__A1 (.I(_1708_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8332__A2 (.I(_2641_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8333__A1 (.I(_2368_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8333__A2 (.I(_1490_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8333__B (.I(_1508_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8333__C (.I(_2651_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8334__A1 (.I(_2494_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8334__A2 (.I(_3424_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8334__B1 (.I(_3433_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8334__B2 (.I(_2352_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8334__C (.I(_3434_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8335__A1 (.I(_2793_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8335__B (.I(_3076_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8336__A1 (.I(_3156_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8336__A2 (.I(_3425_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8339__A1 (.I(_0508_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8339__A2 (.I(_0366_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8340__A1 (.I(_1147_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8340__A2 (.I(_3157_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8341__A1 (.I(_3181_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8341__A2 (.I(_3440_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8341__B (.I(_3441_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8341__C (.I(_2925_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8342__A1 (.I(_2854_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8342__A2 (.I(_3425_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8342__B (.I(_3442_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8342__C (.I(_3058_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8343__A1 (.I(_3293_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8343__A3 (.I(_3443_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8344__A1 (.I(_3415_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8344__A2 (.I(_3424_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8344__B1 (.I(_3433_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8344__B2 (.I(_2524_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8344__C (.I(_2856_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8346__A1 (.I(\as2650.stack[3][3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8346__A2 (.I(_1919_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8346__B1 (.I(_1638_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8347__A1 (.I(\as2650.stack[0][3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8347__C (.I(_0328_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8348__B2 (.I(\as2650.stack[5][3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8349__A2 (.I(_1919_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8349__B1 (.I(_1638_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8349__C (.I(_4475_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8350__A2 (.I(_3448_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8350__B1 (.I(_3449_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8351__A1 (.I(_3426_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8351__A2 (.I(_3425_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8351__B2 (.I(_3446_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8351__C1 (.I(_3451_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8351__C2 (.I(_3327_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8352__A1 (.I(_3371_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8352__B (.I(_3420_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8353__A1 (.I(_3333_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8353__A2 (.I(_3425_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8354__A1 (.I(_0928_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8354__A2 (.I(_3289_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8354__C (.I(_3112_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8355__A2 (.I(_3423_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8356__A1 (.I(_2188_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8356__A2 (.I(_3455_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8357__I (.I(_3456_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8358__I (.I(_3393_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8359__I (.I(_3394_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8360__A2 (.I(_3428_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8361__A2 (.I(_3428_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8362__B (.I(_1685_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8363__A1 (.I(_2188_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8363__A2 (.I(_1605_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8364__A1 (.I(_1679_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8364__A2 (.I(_2698_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8365__A1 (.I(_3256_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8365__A2 (.I(_3457_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8365__B1 (.I(_3464_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8365__B2 (.I(_2524_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8365__C (.I(_2927_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8366__A1 (.I(_0506_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8366__A2 (.I(_0366_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8367__A1 (.I(_0506_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8367__A2 (.I(_0366_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8369__A1 (.I(_1581_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8369__A2 (.I(_0496_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8369__A3 (.I(_3468_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8370__A1 (.I(_0596_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8370__A2 (.I(_1490_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8371__A1 (.I(_1267_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8371__A2 (.I(_0898_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8372__A1 (.I(_2648_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8372__A2 (.I(_3469_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8372__B (.I(_3470_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8372__C (.I(_3471_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8373__A1 (.I(_2353_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8373__A2 (.I(_3464_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8374__A1 (.I(\as2650.addr_buff[4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8374__A2 (.I(_2754_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8375__A1 (.I(_1582_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8375__A2 (.I(_2533_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8375__B (.I(_1508_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8376__A1 (.I(_3082_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8376__A2 (.I(_3456_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8376__B (.I(_3475_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8377__A1 (.I(_2482_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8377__A2 (.I(_2354_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8378__A1 (.I(_3472_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8379__A1 (.I(_3459_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8380__A1 (.I(_3458_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8380__A2 (.I(_3457_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8380__B2 (.I(_3291_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8381__I (.I(_2391_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8382__A1 (.I(\as2650.stack[3][4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8382__A2 (.I(_2215_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8382__B (.I(_4473_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8383__A2 (.I(_1639_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8384__A2 (.I(_1904_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8384__B1 (.I(_1656_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8385__A2 (.I(_3319_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8385__B1 (.I(_3322_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8385__C2 (.I(\as2650.stack[5][4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8386__A1 (.I(_0525_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8387__A1 (.I(\as2650.stack[7][4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8387__A2 (.I(_1920_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8389__A1 (.I(_3481_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8389__A2 (.I(_3488_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8391__A1 (.I(_3210_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8391__A2 (.I(_3457_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8392__I (.I(_2388_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8393__A1 (.I(_3492_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8393__A2 (.I(_3457_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8393__B (.I(_3288_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8394__A1 (.I(_0933_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8394__A2 (.I(_3374_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8394__C (.I(_2415_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8395__A1 (.I(_0933_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8395__A3 (.I(_3423_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8397__I (.I(_3495_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8398__A1 (.I(_3393_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8399__A1 (.I(_1579_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8399__A2 (.I(_2762_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8400__A1 (.I(_0939_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8400__A2 (.I(_1614_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8401__A1 (.I(_4265_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8401__A2 (.I(_3157_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8402__A1 (.I(_0685_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8402__A2 (.I(_2539_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8402__B (.I(_2396_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8403__A1 (.I(_2996_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8403__B1 (.I(_3500_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8404__A1 (.I(_3221_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8404__A2 (.I(_3499_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8404__C (.I(_1294_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8405__I (.I(_3471_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8406__A1 (.I(_2694_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8406__A2 (.I(_0496_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8407__A1 (.I(_2694_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8407__A2 (.I(_0496_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8408__A2 (.I(_3468_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8409__A1 (.I(_1180_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8409__A2 (.I(_0583_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8410__A1 (.I(_2509_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8410__A2 (.I(_3508_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8411__A1 (.I(_2736_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8411__A2 (.I(_2756_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8411__B (.I(_3504_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8411__C (.I(_3509_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8412__A1 (.I(_2196_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8412__A3 (.I(_3428_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8413__A1 (.I(_0940_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8414__A1 (.I(_3395_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8415__A1 (.I(_3059_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8415__B (.I(_3510_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8415__C (.I(_3513_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8416__B (.I(_3391_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8417__A1 (.I(_3250_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8417__A2 (.I(_3495_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8417__B1 (.I(_3499_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8417__B2 (.I(_2513_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8417__C (.I(_3154_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8420__A1 (.I(\as2650.stack[3][5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8420__A2 (.I(_2215_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8421__A2 (.I(_3361_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8421__B1 (.I(_3362_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8421__B2 (.I(\as2650.stack[1][5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8422__A2 (.I(_0426_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8422__B2 (.I(_4453_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8423__A2 (.I(_3366_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8423__B1 (.I(_3386_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8424__A2 (.I(_1904_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8424__B1 (.I(_1656_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8424__B2 (.I(\as2650.stack[5][5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8425__A1 (.I(_0525_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8426__A2 (.I(_3524_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8427__I (.I(_3290_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8428__A1 (.I(_3336_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8428__B1 (.I(_3525_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8428__B2 (.I(_3369_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8428__C (.I(_3526_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8429__A1 (.I(_3379_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8429__A2 (.I(_3495_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8429__C (.I(_3373_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8430__A1 (.I(_0940_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8430__A2 (.I(_3289_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8430__C (.I(_3112_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8432__A1 (.I(_0946_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8432__A2 (.I(_3529_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8433__A1 (.I(_0946_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8433__A2 (.I(_1618_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8434__A1 (.I(_1709_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8434__A2 (.I(_2790_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8435__I (.I(_2645_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8436__A1 (.I(_0759_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8436__A2 (.I(_2539_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8437__A1 (.I(_4357_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8437__A2 (.I(_3345_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8438__A1 (.I(_2495_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8438__B2 (.I(_3533_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8438__C1 (.I(_3089_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8438__C2 (.I(_3535_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8439__A1 (.I(_0758_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8439__A2 (.I(_0674_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8440__A1 (.I(_2800_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8440__A2 (.I(_0583_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8441__A1 (.I(_2800_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8441__A2 (.I(_0583_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8444__B (.I(_3181_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8445__A1 (.I(_1526_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8445__A2 (.I(_2777_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8445__B1 (.I(_3541_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8445__B2 (.I(_3542_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8445__C (.I(_3070_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8446__A1 (.I(_3164_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8446__B (.I(_3543_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8447__A1 (.I(_0946_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8448__A1 (.I(_3459_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8449__A1 (.I(_3458_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8449__B2 (.I(_3126_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8449__C (.I(_3546_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8450__A1 (.I(_3250_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8450__B2 (.I(_2513_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8450__C (.I(_3154_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8451__A1 (.I(_3153_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8452__A1 (.I(_0947_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8452__A2 (.I(_3529_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8453__A2 (.I(_3319_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8455__A2 (.I(_1920_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8455__B1 (.I(_3386_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8456__A2 (.I(_3366_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8456__B1 (.I(_3386_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8457__A1 (.I(\as2650.stack[4][6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8457__A2 (.I(_1904_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8457__B1 (.I(_1656_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8457__B2 (.I(\as2650.stack[5][6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8457__C (.I(_4476_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8458__A1 (.I(_4477_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8460__A1 (.I(_3216_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8460__B1 (.I(_3557_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8460__B2 (.I(_3481_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8460__C (.I(_3371_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8461__A1 (.I(_3333_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8461__C (.I(_3288_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8462__A1 (.I(_2201_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8462__A2 (.I(_3377_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8462__B (.I(_1566_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8463__A2 (.I(_3560_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8464__A1 (.I(_0945_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8464__A2 (.I(_2194_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8465__A1 (.I(_0953_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8465__A2 (.I(_3561_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8466__I (.I(_3562_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8467__A1 (.I(_2825_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8467__A2 (.I(_0674_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8468__A1 (.I(_2825_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8468__A2 (.I(_0674_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8470__A1 (.I(_1604_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8470__A2 (.I(_4370_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8470__A3 (.I(_3566_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8471__A1 (.I(_3345_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8472__A1 (.I(_1619_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8472__A2 (.I(_2540_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8472__B (.I(_3504_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8472__C (.I(_3568_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8473__A1 (.I(_0945_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8473__A3 (.I(_2187_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8474__A1 (.I(_2203_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8474__A2 (.I(_3570_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8475__A1 (.I(_2925_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8475__A2 (.I(_3163_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8475__B (.I(_3156_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8476__A1 (.I(_0953_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8476__A2 (.I(_1605_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8477__A1 (.I(_1679_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8477__A2 (.I(_2849_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8478__A1 (.I(_2153_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8478__A2 (.I(_1489_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8479__A1 (.I(_1599_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8479__A2 (.I(_1490_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8480__A1 (.I(_2526_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8480__A2 (.I(_3562_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8480__B1 (.I(_3576_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8480__B2 (.I(_1509_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8480__C (.I(_2481_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8481__A1 (.I(_2645_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8481__A2 (.I(_3574_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8481__B (.I(_3577_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8481__C (.I(_3076_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8482__A1 (.I(_3395_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8482__B2 (.I(_3572_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8483__A1 (.I(_3293_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8483__A2 (.I(_3569_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8484__A1 (.I(_3415_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8485__A1 (.I(_2492_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8485__A2 (.I(_3574_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8485__C (.I(_3001_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8486__A1 (.I(\as2650.stack[3][7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8486__A2 (.I(_1920_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8486__B1 (.I(_1639_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8487__A2 (.I(_1905_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8487__B1 (.I(_1657_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8487__B2 (.I(\as2650.stack[1][7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8487__C (.I(_0525_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8488__A1 (.I(\as2650.stack[7][7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8488__A2 (.I(_3366_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8488__B1 (.I(_3361_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8488__C1 (.I(\as2650.stack[5][7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8488__C2 (.I(_3362_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8490__A2 (.I(_1639_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8490__B (.I(_4476_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8492__A1 (.I(_3317_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8492__C1 (.I(_3588_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8492__C2 (.I(_2391_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8493__A1 (.I(_3371_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8493__B (.I(_3376_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8494__A1 (.I(_3333_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8495__I (.I(_2577_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8496__A1 (.I(_0953_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8496__A2 (.I(_3289_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8496__C (.I(_3592_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8497__A1 (.I(_0966_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8497__A2 (.I(_3374_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8498__A2 (.I(_3561_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8499__A2 (.I(_3594_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8501__A1 (.I(\as2650.pc[8] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8501__A2 (.I(_2203_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8501__A3 (.I(_3570_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8503__A1 (.I(_2204_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8503__A2 (.I(_3570_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8504__A1 (.I(_3103_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8504__A2 (.I(_3598_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8504__A3 (.I(_3353_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8505__A2 (.I(_1618_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8506__A1 (.I(_1709_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8506__A2 (.I(_2903_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8507__A1 (.I(_1549_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8507__A2 (.I(_2539_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8508__A1 (.I(_2334_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8508__A2 (.I(_2755_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8508__B (.I(_1509_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8509__A1 (.I(_2996_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8510__A1 (.I(_3533_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8510__B (.I(_3604_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8511__A2 (.I(_4370_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8512__A2 (.I(_4370_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8513__A2 (.I(_3566_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8514__A1 (.I(_0896_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8515__A1 (.I(_2899_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8515__A2 (.I(_3610_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8516__A1 (.I(_3598_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8516__B1 (.I(_3611_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8516__B2 (.I(_3070_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8517__B1 (.I(_3596_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8517__B2 (.I(_3572_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8517__C1 (.I(_1443_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8518__A1 (.I(_3257_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8518__A2 (.I(_3596_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8518__B2 (.I(_2550_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8518__C (.I(_2928_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8519__A1 (.I(_3391_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8520__A1 (.I(_3426_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8520__A2 (.I(_3596_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8521__A1 (.I(_1085_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8521__A2 (.I(_1499_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8521__B (.I(_3046_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8522__A1 (.I(_3210_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8522__A2 (.I(_3596_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8522__C (.I(_3420_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8523__I (.I(_1391_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8524__B (.I(_3619_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8526__I (.I(_3288_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8527__A2 (.I(_3594_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8529__I (.I(_3623_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8530__A1 (.I(_2382_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8530__A2 (.I(_3058_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8531__A2 (.I(_3610_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8532__A1 (.I(_2362_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8534__A1 (.I(_0979_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8534__A2 (.I(_1708_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8535__A1 (.I(_1336_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8536__A1 (.I(_3221_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8537__A1 (.I(\as2650.addr_buff[1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8537__A2 (.I(_2538_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8538__A1 (.I(_1275_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8538__A3 (.I(_3632_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8539__A1 (.I(_2526_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8539__A2 (.I(_3623_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8539__B (.I(_3633_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8539__C (.I(_1234_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8540__A1 (.I(_3076_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8540__A3 (.I(_3634_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8540__B (.I(_3095_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8541__A1 (.I(_3572_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8541__A2 (.I(_3624_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8541__B2 (.I(_3395_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8542__A1 (.I(_3625_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8542__A2 (.I(_3627_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8543__A1 (.I(_3257_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8543__A2 (.I(_3624_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8543__B2 (.I(_2549_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8543__C (.I(_2928_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8546__A1 (.I(_0335_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8546__A2 (.I(_3369_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8546__B1 (.I(_3317_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8546__B2 (.I(_3624_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8547__B (.I(_3329_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8548__A1 (.I(_3292_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8548__A2 (.I(_3624_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8548__C (.I(_3331_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8549__A2 (.I(_3621_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8549__C (.I(_3592_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8550__A2 (.I(\as2650.pc[8] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8550__A3 (.I(_3594_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8551__A1 (.I(_2969_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8551__A2 (.I(_3644_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8552__A1 (.I(_2952_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8552__A2 (.I(_3610_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8553__A1 (.I(_2365_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8555__A1 (.I(_2969_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8555__A2 (.I(_3648_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8556__A1 (.I(_0990_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8556__A2 (.I(_1544_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8557__A1 (.I(_1709_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8557__A2 (.I(_2976_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8558__A1 (.I(_0989_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8558__A2 (.I(_3644_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8559__A1 (.I(_2395_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8559__A2 (.I(_3406_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8560__A1 (.I(_2365_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8560__A2 (.I(_2776_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8561__A1 (.I(_2527_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8561__A2 (.I(_3652_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8561__B (.I(_3654_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8561__C (.I(_2160_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8562__A1 (.I(_3533_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8563__A1 (.I(_3504_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8563__A2 (.I(_3647_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8563__B2 (.I(_3459_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8563__C1 (.I(_3103_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8564__A1 (.I(_3458_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8564__C (.I(_3391_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8565__A1 (.I(_3250_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8565__B2 (.I(_2492_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8565__C (.I(_3001_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8567__A1 (.I(_0436_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8567__A2 (.I(_3481_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8567__B1 (.I(_3426_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8567__B2 (.I(_3652_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8567__C (.I(_3526_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8568__A1 (.I(_3379_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8568__B2 (.I(_3661_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8568__C (.I(_3373_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8569__A1 (.I(_2969_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8569__A2 (.I(_3621_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8569__B (.I(_3662_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8569__C (.I(_3592_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8570__A2 (.I(_3644_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8571__A2 (.I(_3663_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8573__A1 (.I(_0989_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8573__A2 (.I(_3648_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8575__A1 (.I(_2950_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8575__A2 (.I(_3610_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8575__B (.I(_2369_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8576__A1 (.I(_2998_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8576__A2 (.I(_2538_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8576__A3 (.I(_3021_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8577__A2 (.I(_3669_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8578__A1 (.I(_3392_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8578__A2 (.I(_3665_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8579__A1 (.I(_3459_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8579__B1 (.I(_3670_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8579__B2 (.I(_3504_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8580__I1 (.I(_3006_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8580__S (.I(_0837_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8581__A1 (.I(_3533_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8582__A1 (.I(_2368_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8582__A2 (.I(_2385_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8582__B (.I(_3441_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8583__A1 (.I(_2481_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8583__A2 (.I(_2354_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8584__A1 (.I(_2495_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8584__A2 (.I(_3665_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8584__B1 (.I(_3675_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8584__B2 (.I(_1277_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8584__C (.I(_3676_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8585__A1 (.I(_3256_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8585__B2 (.I(_2524_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8585__C (.I(_2927_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8587__A1 (.I(_3153_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8588__A1 (.I(_0533_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8588__A2 (.I(_3327_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8588__B1 (.I(_3317_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8588__B2 (.I(_3665_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8589__B (.I(_3526_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8590__A1 (.I(_3292_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8590__A2 (.I(_3665_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8590__C (.I(_3331_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8591__A1 (.I(_2995_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8591__A2 (.I(_3621_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8591__C (.I(_3592_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8592__A1 (.I(\as2650.pc[11] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8592__A2 (.I(_3663_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8593__A1 (.I(_3035_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8595__A1 (.I(_0995_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8595__A3 (.I(_3648_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8596__A1 (.I(_1003_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8596__A2 (.I(_3687_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8597__A1 (.I(_3020_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8597__A2 (.I(_3669_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8598__A1 (.I(_3394_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8598__B1 (.I(_3689_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8598__B2 (.I(_3471_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8599__I1 (.I(_3017_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8599__S (.I(_1599_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8600__A1 (.I(_2353_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8601__A1 (.I(_2372_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8601__A2 (.I(_2776_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8601__B (.I(_3470_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8602__A1 (.I(_3082_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8602__A2 (.I(_3686_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8602__B1 (.I(_3693_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8602__B2 (.I(_1276_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8602__C (.I(_3676_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8603__A1 (.I(_3256_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8603__B2 (.I(_2523_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8603__C (.I(_2855_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8605__A1 (.I(_3194_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8606__A1 (.I(_3046_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8607__A1 (.I(_3458_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8607__A2 (.I(_3686_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8608__A1 (.I(_0632_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8608__A2 (.I(_1499_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8609__A1 (.I(_3210_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8609__A2 (.I(_3686_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8610__A1 (.I(_3492_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8610__A2 (.I(_3686_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8610__B (.I(_3331_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8611__A1 (.I(_3035_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8611__A2 (.I(_3374_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8611__C (.I(_2415_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8612__I (.I(_2415_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8613__A2 (.I(_0995_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8613__A3 (.I(_3663_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8615__I (.I(_3705_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8616__A1 (.I(_3035_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8616__A2 (.I(_3687_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8618__I1 (.I(_3705_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8618__S (.I(_3353_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8619__A1 (.I(_1251_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8619__A2 (.I(_3709_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8620__A1 (.I(_2996_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8620__A2 (.I(_3705_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8621__A1 (.I(_1008_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8621__A2 (.I(_1544_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8622__A1 (.I(_4265_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8622__A2 (.I(_3345_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8622__B1 (.I(_2353_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8622__B2 (.I(_3712_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8622__C (.I(_3048_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8623__A3 (.I(_3713_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8624__A1 (.I(_3093_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8625__A1 (.I(_2372_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8625__A2 (.I(_3669_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8625__B (.I(_3500_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8625__C (.I(_2382_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8626__A1 (.I(_2926_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8626__A2 (.I(_3706_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8626__C (.I(_3598_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8627__A1 (.I(_3257_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8627__A2 (.I(_3706_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8627__B1 (.I(_3712_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8627__B2 (.I(_2549_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8627__C (.I(_2856_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8629__A1 (.I(_0709_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8629__A2 (.I(_3481_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8629__B1 (.I(_3426_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8629__B2 (.I(_3706_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8630__A1 (.I(_3329_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8630__A2 (.I(_3706_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8631__A1 (.I(_3379_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8631__C (.I(_3420_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8632__A1 (.I(_1008_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8632__A2 (.I(_3377_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8633__A1 (.I(_3703_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8634__I (.I(\as2650.pc[14] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8635__A3 (.I(_0995_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8635__A4 (.I(_3663_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8636__A1 (.I(_3724_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8638__A1 (.I(_4264_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8638__A2 (.I(_3158_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8638__B (.I(_3625_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8639__A1 (.I(_1008_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8640__A1 (.I(\as2650.pc[14] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8641__I (.I(_3081_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8642__A1 (.I(_4264_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8642__A2 (.I(_2410_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8642__B1 (.I(_2494_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8642__C2 (.I(\as2650.pc[14] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8643__B2 (.I(_2482_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8644__A1 (.I(_3393_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8644__A2 (.I(_3727_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8644__B1 (.I(_3733_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8644__B2 (.I(_3598_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8645__B (.I(_3293_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8646__A1 (.I(_2634_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8646__A2 (.I(_3727_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8647__A1 (.I(_3724_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8647__A2 (.I(_3148_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8647__C (.I(_3194_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8648__A1 (.I(_3214_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8649__A1 (.I(_0781_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8649__A2 (.I(_3327_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8649__B1 (.I(_2388_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8649__B2 (.I(_3727_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8650__B (.I(_3526_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8651__A1 (.I(_3292_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8651__A2 (.I(_3727_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8651__C (.I(_3373_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8652__I (.I(_2577_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8653__A1 (.I(_3724_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8653__A2 (.I(_3621_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8653__C (.I(_3742_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8654__A1 (.I(_1453_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8654__A2 (.I(_2420_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8655__A1 (.I(_1329_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8655__A2 (.I(_2472_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8655__B (.I(_3265_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8656__A1 (.I(_2755_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8656__A2 (.I(_0600_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8656__B2 (.I(_3175_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8656__C (.I(_4260_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8657__B (.I(_1516_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8658__A1 (.I(_4160_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8658__A2 (.I(_3265_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8658__A3 (.I(_1288_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8659__A1 (.I(_2927_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8659__A2 (.I(_3747_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8659__B (.I(_0971_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8660__A1 (.I(_4419_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8660__A2 (.I(_1046_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8660__B (.I(_4395_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8661__A1 (.I(_1463_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8661__A2 (.I(_3748_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8661__B2 (.I(_3265_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8662__A1 (.I(_1328_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8662__A2 (.I(_1338_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8662__B (.I(_1496_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8662__C (.I(_2448_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8663__A1 (.I(_4242_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8663__A2 (.I(_2469_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8663__A3 (.I(_1491_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8663__B (.I(_3751_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8665__A1 (.I(_1939_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8665__A2 (.I(_0871_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8665__A3 (.I(_1352_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8665__A4 (.I(_1487_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8666__A1 (.I(_1333_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8666__A2 (.I(_1474_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8667__A1 (.I(_1318_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8667__A2 (.I(_1476_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8667__A4 (.I(_1484_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8668__A2 (.I(_3750_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8668__A3 (.I(_3755_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8668__A4 (.I(_3756_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8669__I (.I(_3757_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8670__A1 (.I(_2598_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8670__A2 (.I(_4361_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8671__A1 (.I(_2477_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8671__A2 (.I(_4353_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8672__A1 (.I(_3143_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8672__A2 (.I(_1100_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8672__B (.I(_3080_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8673__A1 (.I(_3219_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8673__A2 (.I(_4344_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8673__B1 (.I(_3183_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8673__B2 (.I(_3760_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8674__I (.I(_3757_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8675__A1 (.I(_4398_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8675__A2 (.I(_2632_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8676__I (.I(_4394_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8677__I (.I(_3765_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8678__I (.I(_1535_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8679__A2 (.I(_3326_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8680__I (.I(_1235_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8681__A1 (.I(_4428_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8682__A1 (.I(_0550_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8682__A2 (.I(_3770_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8682__A3 (.I(_0340_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8685__A1 (.I(_1589_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8685__A2 (.I(_3773_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8686__A1 (.I(_4316_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8686__A2 (.I(_3772_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8687__A1 (.I(_1736_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8687__A2 (.I(_3769_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8687__B1 (.I(_4435_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8688__I (.I(_4219_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8689__A1 (.I(_3768_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8689__B (.I(_3777_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8690__A1 (.I(_1624_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8690__A2 (.I(_4377_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8690__B (.I(_3778_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8690__C (.I(_1535_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8691__I (.I(_4394_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8692__A1 (.I(_3767_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8692__A2 (.I(_1383_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8692__B (.I(_3779_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8692__C (.I(_3780_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8693__A1 (.I(_1691_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8693__A2 (.I(_3766_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8693__B (.I(_2629_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8694__A2 (.I(_3763_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8694__A4 (.I(_3782_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8695__A1 (.I(_4441_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8696__A1 (.I(_3703_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8697__I (.I(_2337_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8698__I0 (.I(_4513_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8698__I1 (.I(_0292_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8699__A1 (.I(_3143_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8699__A2 (.I(_1383_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8699__B (.I(_3080_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8700__A1 (.I(_3219_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8700__A2 (.I(_0321_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8700__B1 (.I(_3183_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8700__B2 (.I(_3786_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8701__A1 (.I(_1552_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8701__A2 (.I(_1541_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8701__B (.I(_3170_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8702__I (.I(_4227_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8703__A2 (.I(_3368_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8704__I (.I(_2423_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8705__I (.I(_3792_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8706__A1 (.I(\as2650.psl[1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8706__A2 (.I(_3792_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8707__A1 (.I(_4458_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8707__A2 (.I(_3793_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8708__A1 (.I(_1733_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8708__A2 (.I(_3769_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8708__B1 (.I(_4435_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8708__C (.I(_3777_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8709__A1 (.I(_1519_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8709__A2 (.I(_4514_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8709__B (.I(_1480_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8710__A1 (.I(_3791_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8710__A2 (.I(_3796_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8710__B (.I(_3797_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8711__A2 (.I(_0400_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8711__B (.I(_3798_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8711__C (.I(_3765_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8712__A1 (.I(_3199_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8712__A2 (.I(_4535_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8713__A1 (.I(_3088_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8714__A1 (.I(_3763_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8714__A2 (.I(_3788_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8715__A1 (.I(_1382_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8716__A1 (.I(_3703_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8717__I (.I(_2337_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8718__A2 (.I(_0358_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8719__A1 (.I(_3804_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8719__A2 (.I(_2592_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8720__A1 (.I(_3143_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8720__A2 (.I(_4527_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8720__B (.I(_3080_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8721__A1 (.I(_3219_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8721__A2 (.I(_0422_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8721__B1 (.I(_3183_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8721__B2 (.I(_3806_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8722__A1 (.I(_0378_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8722__A2 (.I(_2632_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8723__I (.I(_1623_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8724__A2 (.I(_3390_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8726__A1 (.I(_0849_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8726__A2 (.I(_3773_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8727__A1 (.I(_3812_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8727__A2 (.I(_3772_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8728__A1 (.I(_3769_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8728__A2 (.I(_1749_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8728__B2 (.I(_4435_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8728__C (.I(_1623_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8729__A1 (.I(_3810_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8729__A2 (.I(_4388_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8729__B1 (.I(_3811_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8729__B2 (.I(_3815_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8731__A1 (.I(_3767_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8731__A2 (.I(_1393_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8731__B (.I(_3817_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8731__C (.I(_3765_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8732__A1 (.I(_1699_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8732__A2 (.I(_3766_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8732__B (.I(_2629_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8733__A1 (.I(_3763_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8734__A1 (.I(_0917_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8735__A1 (.I(_3703_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8736__A1 (.I(_2338_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8736__A2 (.I(_0491_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8737__A2 (.I(_0485_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8737__C (.I(_2756_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8738__A1 (.I(_2756_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8738__A2 (.I(_0476_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8738__C (.I(_3126_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8739__A1 (.I(_3144_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8739__A2 (.I(_1393_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8739__B (.I(_3824_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8739__C (.I(_3088_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8740__A2 (.I(_3451_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8741__I (.I(_4365_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8742__A1 (.I(\as2650.psu[3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8743__A1 (.I(_3827_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8743__A2 (.I(_3773_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8744__A1 (.I(_1235_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8744__A2 (.I(_1764_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8744__B2 (.I(_4434_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8745__A1 (.I(_3826_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8745__B (.I(_3777_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8746__A1 (.I(_3810_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8746__A2 (.I(_0400_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8746__B (.I(_3831_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8746__C (.I(_1535_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8747__A2 (.I(_0694_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8747__C (.I(_3765_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8748__A1 (.I(_1556_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8748__A2 (.I(_3780_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8748__B (.I(_2629_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8748__C (.I(_3833_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8749__A1 (.I(_0512_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8749__A2 (.I(_2753_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8749__B (.I(_3757_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8749__C (.I(_3834_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8750__A1 (.I(_0924_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8751__A1 (.I(_3189_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8751__A2 (.I(_3836_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8752__I (.I(_3763_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8753__I (.I(_2386_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8754__A1 (.I(_3804_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8754__A2 (.I(_0614_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8755__A1 (.I(_2477_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8755__A2 (.I(_0578_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8756__A1 (.I(_1572_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8756__A2 (.I(_0566_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8756__B (.I(_1518_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8757__A1 (.I(_3838_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8757__A2 (.I(_0570_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8757__B1 (.I(_3184_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8758__A2 (.I(_3488_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8759__I (.I(_1235_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8760__A1 (.I(\as2650.psu[4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8760__A2 (.I(_3772_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8761__A1 (.I(_1033_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8761__A2 (.I(_3772_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8762__I (.I(_4434_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8763__A1 (.I(_3844_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8763__A2 (.I(_2027_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8763__B1 (.I(_3846_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8763__B2 (.I(_3847_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8763__C (.I(_3810_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8764__A1 (.I(_1520_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8764__A2 (.I(_0372_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8765__A1 (.I(_3843_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8765__A2 (.I(_3848_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8765__C (.I(_3767_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8766__I (.I(_1628_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8767__A1 (.I(_3851_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8767__A2 (.I(_0593_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8767__B (.I(_1541_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8768__A1 (.I(_1558_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8768__A2 (.I(_1547_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8768__B1 (.I(_3850_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8768__B2 (.I(_3852_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8768__C (.I(_1513_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8769__A1 (.I(_0603_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8769__A2 (.I(_2633_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8770__A1 (.I(_3842_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8771__I (.I(_3757_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8772__A1 (.I(_0579_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8772__A2 (.I(_3856_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8772__B (.I(_3245_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8773__A1 (.I(_3837_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8774__A1 (.I(_2598_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8774__A2 (.I(_0698_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8775__A1 (.I(_3804_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8775__A2 (.I(_0668_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8776__A1 (.I(_2399_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8776__A2 (.I(_0639_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8776__B (.I(_2514_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8777__A1 (.I(_3838_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8777__A2 (.I(_0662_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8777__B1 (.I(_3184_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8778__A1 (.I(_3810_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8778__A2 (.I(_0694_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8779__A1 (.I(\as2650.psl[5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8779__A2 (.I(_3792_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8780__A1 (.I(_1226_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8780__A2 (.I(_3793_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8781__A1 (.I(_3769_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8781__A2 (.I(_1812_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8781__B2 (.I(_3847_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8781__C (.I(_1623_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8782__A1 (.I(_0341_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8782__A2 (.I(_3525_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8782__B (.I(_3865_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8783__A2 (.I(_3866_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8784__A1 (.I(_1628_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8784__A2 (.I(_1537_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8785__A1 (.I(_3780_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8785__A2 (.I(_3867_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8785__A3 (.I(_3868_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8786__A1 (.I(_1292_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8786__A2 (.I(_3766_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8787__A1 (.I(_0690_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8787__A2 (.I(_2633_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8787__B2 (.I(_2630_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8789__A1 (.I(_0711_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8789__A2 (.I(_3856_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8789__B (.I(_3245_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8790__A1 (.I(_3837_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8790__A2 (.I(_3872_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8791__A1 (.I(_2565_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8791__A2 (.I(_0771_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8792__A1 (.I(_3804_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8792__A2 (.I(_0749_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8793__A1 (.I(_2635_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8793__A2 (.I(_1537_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8793__B (.I(_1450_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8794__A1 (.I(_3838_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8794__A2 (.I(_0740_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8794__B1 (.I(_3184_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8795__I0 (.I(net27));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8795__I1 (.I(_1525_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8795__S (.I(_3792_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8796__A1 (.I(_3844_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8796__A2 (.I(_2084_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8796__B2 (.I(_3847_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8796__C (.I(_3777_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8797__A1 (.I(_0342_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8797__A2 (.I(_3557_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8797__B (.I(_3879_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8798__A1 (.I(_1627_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8798__A2 (.I(_0639_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8798__B (.I(_3880_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8798__C (.I(_3851_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8799__A1 (.I(_3767_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8799__A2 (.I(_0818_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8799__B (.I(_3780_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8800__A1 (.I(_1588_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8800__A2 (.I(_3766_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8800__C (.I(_2630_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8801__A1 (.I(_2458_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8801__A2 (.I(_2753_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8802__A1 (.I(_0944_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8802__A2 (.I(_3856_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8802__B (.I(_3245_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8803__A1 (.I(_3837_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8803__A2 (.I(_3884_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8804__A1 (.I(_2338_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8804__A2 (.I(_0830_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8805__A2 (.I(_0828_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8806__A1 (.I(_2635_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8806__A2 (.I(_0818_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8806__B (.I(_3887_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8806__C (.I(_2514_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8807__A1 (.I(_3838_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8807__A2 (.I(_1212_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8808__A1 (.I(_0620_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8808__A2 (.I(_3588_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8809__A1 (.I(_1611_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8809__A2 (.I(_3793_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8810__A1 (.I(_3262_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8810__A2 (.I(_3793_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8811__A1 (.I(_2109_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8811__A2 (.I(_3844_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8811__B1 (.I(_3847_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8811__C (.I(_1624_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8812__A1 (.I(_3890_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8812__A2 (.I(_3893_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8812__B (.I(_1629_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8813__A2 (.I(_3894_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8814__A1 (.I(_2630_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8814__A2 (.I(_1548_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8814__A3 (.I(_3895_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8815__A1 (.I(_0834_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8815__A2 (.I(_2753_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8816__A1 (.I(_1411_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8816__A2 (.I(_3856_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8816__B (.I(_1634_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8817__A1 (.I(_3837_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8817__A2 (.I(_3897_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8818__A1 (.I(_0957_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8818__A2 (.I(_0427_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8819__A1 (.I(_2208_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8820__I (.I(_3900_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8823__I (.I(_3903_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8824__A1 (.I(_2223_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8824__A2 (.I(_0626_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8824__A3 (.I(_0901_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8825__I (.I(_3905_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8826__A1 (.I(_2146_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8827__A1 (.I(_0848_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8828__I (.I(_3903_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8829__I (.I(_3905_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8830__I (.I(_3900_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8831__A1 (.I(_2285_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8831__A2 (.I(_3908_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8831__B1 (.I(_3909_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8831__C (.I(_3910_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8832__A1 (.I(_2223_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8832__A2 (.I(_0624_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8832__A3 (.I(_0968_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8833__A1 (.I(_2290_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8833__A2 (.I(_3912_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8835__A1 (.I(_2258_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8835__A2 (.I(_3908_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8835__B1 (.I(_3909_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8835__C (.I(_3910_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8836__A1 (.I(_2294_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8836__A2 (.I(_3912_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8838__A1 (.I(_2296_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8838__A2 (.I(_3908_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8838__B1 (.I(_3909_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8838__C (.I(_3910_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8839__A1 (.I(_2298_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8839__A2 (.I(_3912_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8841__A1 (.I(_2300_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8842__A1 (.I(_0932_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8843__A1 (.I(_2302_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8844__A1 (.I(_0938_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8845__A1 (.I(_2265_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8845__C (.I(_3910_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8846__A1 (.I(_2199_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8847__A1 (.I(_2305_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8847__A2 (.I(_3908_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8847__B1 (.I(_3909_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8847__C (.I(_3900_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8848__A1 (.I(_2307_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8848__A2 (.I(_3912_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8851__I (.I(_3923_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8854__I (.I(_3926_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8855__A2 (.I(_0624_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8855__A3 (.I(_0901_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8856__I (.I(_3928_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8857__A1 (.I(_2146_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8857__B2 (.I(\as2650.stack[7][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8858__A1 (.I(_0848_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8859__I (.I(_3926_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8860__I (.I(_3928_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8861__I (.I(_3923_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8862__A1 (.I(_2285_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8862__A2 (.I(_3931_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8862__C (.I(_3933_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8863__A1 (.I(_0968_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8864__A1 (.I(_2290_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8864__A2 (.I(_3935_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8866__A1 (.I(_0921_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8866__A2 (.I(_3931_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8866__C (.I(_3933_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8867__A1 (.I(_2294_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8867__A2 (.I(_3935_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8869__A1 (.I(_2296_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8869__A2 (.I(_3931_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8869__C (.I(_3933_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8870__A1 (.I(_2298_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8870__A2 (.I(_3935_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8872__A1 (.I(_2300_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8872__B2 (.I(\as2650.stack[7][4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8873__A1 (.I(_0932_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8874__A1 (.I(_2302_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8875__A1 (.I(_0938_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8876__A1 (.I(_0948_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8876__C (.I(_3933_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8877__A1 (.I(_2199_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8878__A1 (.I(_2305_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8878__A2 (.I(_3931_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8878__B2 (.I(\as2650.stack[7][7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8878__C (.I(_3923_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8879__A1 (.I(_2307_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8879__A2 (.I(_3935_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8881__A1 (.I(_1019_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8882__I (.I(_3946_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8883__I (.I(_3947_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8884__I (.I(_3947_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8885__A2 (.I(_3949_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8886__A1 (.I(_1653_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8886__A2 (.I(_3948_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8887__I (.I(_3946_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8888__A1 (.I(\as2650.stack[7][9] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8889__A1 (.I(_1663_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8889__A2 (.I(_3948_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8891__A1 (.I(_1666_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8891__A2 (.I(_3948_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8893__A1 (.I(_1668_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8893__A2 (.I(_3948_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8895__A1 (.I(_1670_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8895__A2 (.I(_3949_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8896__A1 (.I(\as2650.stack[7][13] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8896__A2 (.I(_3947_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8897__A1 (.I(_1672_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8897__A2 (.I(_3949_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8898__A2 (.I(_3947_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8899__A1 (.I(_1674_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8899__A2 (.I(_3949_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8900__A1 (.I(_1601_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8900__A2 (.I(_4272_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8901__I (.I(_3958_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8902__A1 (.I(_4153_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8902__A2 (.I(_4491_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8904__I (.I(_3961_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8905__A1 (.I(_1390_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8905__A3 (.I(_3958_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8907__A1 (.I(_3962_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8907__B1 (.I(_3964_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8907__B2 (.I(\as2650.r123[1][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8908__A1 (.I(_4414_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8908__A2 (.I(_3959_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8909__I (.I(_3961_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8911__A1 (.I(_3966_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8911__A2 (.I(_1738_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8911__B1 (.I(_3967_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8912__I (.I(_3958_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8913__A1 (.I(_0323_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8913__A2 (.I(_3969_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8915__A1 (.I(_3966_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8915__A2 (.I(_1753_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8915__B1 (.I(_3967_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8916__A1 (.I(_0424_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8916__A2 (.I(_3969_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8918__A1 (.I(_3962_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8918__A2 (.I(_1772_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8918__B1 (.I(_3964_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8919__A1 (.I(_0523_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8919__A2 (.I(_3959_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8920__A1 (.I(_3962_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8920__B1 (.I(_3964_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8921__A1 (.I(_0616_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8921__A2 (.I(_3969_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8923__A1 (.I(_0981_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8923__A2 (.I(_1939_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8924__A1 (.I(_3976_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8924__A2 (.I(_1823_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8925__A2 (.I(_3967_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8926__A1 (.I(_0703_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8926__A2 (.I(_3969_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8928__A1 (.I(_3976_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8928__A2 (.I(_1859_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8929__A2 (.I(_3967_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8930__A1 (.I(_0775_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8930__A2 (.I(_3958_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8932__A1 (.I(_3976_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8932__A2 (.I(_1898_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8933__A2 (.I(_3964_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8934__A1 (.I(_0846_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8934__A2 (.I(_3959_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8935__A1 (.I(_4272_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8935__A2 (.I(_1612_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8938__A1 (.I(_1390_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8938__A2 (.I(_3961_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8940__A2 (.I(_3989_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8941__A1 (.I(_3966_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8941__A2 (.I(_1979_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8942__A1 (.I(_4414_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8945__A1 (.I(_0323_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8945__A2 (.I(_3992_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8945__B1 (.I(_3993_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8946__I (.I(_3961_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8947__A1 (.I(_3995_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8947__A2 (.I(_2017_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8949__A1 (.I(_0424_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8949__A2 (.I(_3992_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8949__B1 (.I(_3993_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8950__A1 (.I(_3995_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8952__A1 (.I(_0524_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8952__A2 (.I(_3992_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8952__B1 (.I(_3993_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8953__A1 (.I(_3995_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8953__A2 (.I(_2076_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8955__A1 (.I(_0616_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8955__B1 (.I(_3989_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8956__A1 (.I(_3976_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8956__A2 (.I(_2100_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8957__A1 (.I(_0703_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8957__A2 (.I(_3992_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8957__B1 (.I(_3993_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8958__A1 (.I(_3995_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8960__A1 (.I(_0775_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8960__B1 (.I(_3989_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8961__A1 (.I(_3966_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8961__A2 (.I(_2129_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8963__A2 (.I(_3989_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8964__B (.I(_3962_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8965__A1 (.I(_0846_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8965__C (.I(_4007_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8966__A1 (.I(_1556_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8966__A2 (.I(_1704_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8967__A1 (.I(_3191_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8967__A2 (.I(_1698_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8968__A1 (.I(_2373_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8968__A2 (.I(_1704_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8969__A1 (.I(_1570_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8969__A2 (.I(_1698_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8970__A1 (.I(_1555_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8970__A2 (.I(_2634_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8971__A1 (.I(_3191_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8971__A2 (.I(_2509_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8971__A3 (.I(_3048_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8971__A4 (.I(_1309_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8972__A1 (.I(_2926_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8972__A2 (.I(_4011_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8973__A2 (.I(_1481_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8974__A1 (.I(_3045_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8974__C (.I(_3273_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8976__A1 (.I(_1482_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8976__A2 (.I(_3163_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8976__A3 (.I(_0875_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8977__A1 (.I(_1250_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8977__A2 (.I(_3773_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8978__A2 (.I(_1467_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8979__A1 (.I(_1278_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8979__A2 (.I(_1242_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8979__B (.I(_1716_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8979__C (.I(_4018_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8980__A1 (.I(_2342_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8980__A2 (.I(_2400_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8980__A3 (.I(_4016_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8980__A4 (.I(_4019_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8981__A2 (.I(_0897_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8981__B1 (.I(_2408_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8981__B2 (.I(_1272_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8982__A1 (.I(_1498_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8982__A2 (.I(_3236_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8983__A1 (.I(_3844_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8983__A2 (.I(_2449_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8983__A3 (.I(_1281_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8983__A4 (.I(_1357_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8984__A1 (.I(_1046_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8984__A2 (.I(_4020_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8984__A3 (.I(_4022_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8984__A4 (.I(_4023_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8985__A1 (.I(_3415_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8985__A2 (.I(_2438_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8986__A1 (.I(_4012_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8986__A2 (.I(_4015_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8986__A4 (.I(_4025_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8987__A1 (.I(_3336_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8987__A2 (.I(_4010_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8987__B (.I(_4026_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8988__A1 (.I(_2634_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8988__A2 (.I(_3266_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8989__A1 (.I(_0849_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8989__A2 (.I(_0426_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8990__I (.I(_0854_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8991__I0 (.I(_4029_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8991__I1 (.I(_0360_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8992__A1 (.I(_2794_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8992__A2 (.I(_0342_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8993__A1 (.I(_4010_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8993__A2 (.I(_4028_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8994__A1 (.I(_1087_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8994__A2 (.I(_1287_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8995__A1 (.I(_1287_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8995__B2 (.I(_0526_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8995__C (.I(_3199_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8996__A1 (.I(_3230_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8996__A2 (.I(_4029_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8997__A1 (.I(_4027_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8998__A1 (.I(_2223_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8998__A2 (.I(_4027_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__8999__A1 (.I(_3189_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9000__A1 (.I(_3492_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9000__A2 (.I(_3122_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9000__B (.I(_4026_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9001__A1 (.I(_4479_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9001__A2 (.I(_0624_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9002__I (.I(_3122_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9003__A1 (.I(_1921_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9003__A2 (.I(_1640_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9004__A1 (.I(_4042_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9004__B1 (.I(_1009_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9004__B2 (.I(_3123_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9005__A1 (.I(_2635_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9005__A2 (.I(_3266_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9005__B (.I(_4041_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9005__C (.I(_4043_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9006__A1 (.I(_4040_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9006__B1 (.I(_4044_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9006__B2 (.I(_1287_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9006__C (.I(_3230_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9007__A1 (.I(_3230_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9007__A2 (.I(_4040_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9008__A1 (.I(_4463_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9008__B (.I(_1634_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9010__A1 (.I(_3214_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9010__A2 (.I(_1551_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9010__A3 (.I(_3126_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9010__A4 (.I(_1249_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9011__A1 (.I(_4026_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9011__A2 (.I(_4048_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9012__A1 (.I(_0620_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9013__A1 (.I(_4050_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9013__A2 (.I(_3113_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9013__B1 (.I(_3114_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9014__A1 (.I(_0621_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9014__A3 (.I(_3216_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9015__A1 (.I(_3136_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9015__A2 (.I(_3216_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9015__B (.I(_1589_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9016__A1 (.I(_3492_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9016__A2 (.I(_4051_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9017__A1 (.I(_1589_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9018__C (.I(_3742_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9019__A1 (.I(_1517_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9019__A2 (.I(_1622_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9019__A3 (.I(_1624_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9020__A1 (.I(_0553_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9020__A2 (.I(_1364_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9021__A1 (.I(_4491_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9021__A2 (.I(_3268_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9022__A1 (.I(_2776_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9022__A2 (.I(_1317_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9022__C (.I(_4058_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9023__A1 (.I(_1359_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9023__A2 (.I(_4059_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9024__A1 (.I(_1234_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9024__A2 (.I(_1233_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9024__A3 (.I(_1466_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9025__A1 (.I(_2395_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9025__A2 (.I(_1264_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9026__A1 (.I(_1463_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9026__A3 (.I(_4062_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9027__A1 (.I(_1475_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9027__A3 (.I(_4060_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9028__A1 (.I(_0855_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9029__A1 (.I(_4365_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9029__A2 (.I(_1251_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9030__A1 (.I(_3827_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9030__A2 (.I(_0516_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9030__B (.I(_2631_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9030__C (.I(_1034_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9031__A1 (.I(_2450_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9031__A2 (.I(_3074_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9031__A3 (.I(_4067_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9032__A1 (.I(_1163_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9033__A1 (.I(_1476_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9033__A2 (.I(_4064_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9033__A3 (.I(_4065_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9034__A1 (.I(_1291_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9034__A2 (.I(_4056_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9034__B (.I(_4070_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9035__A1 (.I(_4430_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9035__A2 (.I(_1527_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9036__A1 (.I(_4072_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9036__A2 (.I(_1290_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9036__B (.I(_1520_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9037__A1 (.I(_1627_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9037__A2 (.I(_0566_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9037__B1 (.I(_3141_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9038__A1 (.I(_3851_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9038__B (.I(_3868_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9039__A1 (.I(_3088_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9039__A2 (.I(_0570_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9040__A1 (.I(_1451_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9041__C (.I(_3742_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9042__A1 (.I(_1691_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9042__A2 (.I(_4056_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9042__B (.I(_4070_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9044__A2 (.I(_0319_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9046__A1 (.I(_0421_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9046__A2 (.I(_0451_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9046__B1 (.I(_4079_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9046__B2 (.I(_4081_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9047__A1 (.I(_0421_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9047__A2 (.I(_0451_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9047__B1 (.I(_0467_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9048__A1 (.I(_0561_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9048__A2 (.I(_0569_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9049__A1 (.I(_0467_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9049__A2 (.I(_0476_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9050__A1 (.I(_0561_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9050__A2 (.I(_0569_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9050__B1 (.I(_0653_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9050__B2 (.I(_0661_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9051__A1 (.I(_0653_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9051__A2 (.I(_0661_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9051__B1 (.I(_0732_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9052__A1 (.I(_0732_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9053__A1 (.I(_0821_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9053__A2 (.I(_1431_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9054__A1 (.I(_0821_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9054__A2 (.I(_1431_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9054__B (.I(_1518_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9055__A1 (.I(_4072_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9055__A2 (.I(_3113_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9055__B (.I(_1519_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9056__A1 (.I(_1627_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9056__A2 (.I(_0818_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9056__B1 (.I(_3115_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9056__C (.I(_1628_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9057__A1 (.I(_3851_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9057__A2 (.I(_1100_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9058__A1 (.I(_4089_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9058__B1 (.I(_4093_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9058__B2 (.I(_1576_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9059__A1 (.I(_4316_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9059__C (.I(_3742_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9060__A1 (.I(_3106_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9060__A2 (.I(_1046_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9060__A3 (.I(_1244_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9060__A4 (.I(_2631_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9061__A1 (.I(_1575_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9061__A2 (.I(_4010_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9062__A1 (.I(_4064_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9063__A1 (.I(_1212_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9063__A2 (.I(_1431_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9064__A1 (.I(_1518_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9064__A2 (.I(_0801_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9065__I (.I(_4072_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9066__A1 (.I(_4100_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9067__B2 (.I(_1576_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9067__C (.I(_4097_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9068__A1 (.I(_3812_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9068__A2 (.I(_4097_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9068__C (.I(_3249_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9069__A1 (.I(_2793_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9069__A2 (.I(_1469_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9070__A1 (.I(_3770_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9070__A2 (.I(_3268_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9070__A3 (.I(_4062_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9071__A1 (.I(_1270_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9072__A1 (.I(_2373_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9072__A2 (.I(_3144_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9072__B (.I(_4105_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9073__A1 (.I(_1089_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9073__A2 (.I(_4106_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9074__I (.I(_4105_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9075__A1 (.I(_4100_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9076__A1 (.I(_3138_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9077__A2 (.I(_4110_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9077__B (.I(_3619_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9078__A1 (.I(_3132_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9078__A2 (.I(_4105_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9079__A1 (.I(_4365_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9080__I (.I(_1622_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9081__A1 (.I(_4113_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9081__A2 (.I(_4100_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9081__B (.I(_3133_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9083__B (.I(_3619_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9084__A1 (.I(_1552_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9084__A2 (.I(_3136_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9084__A3 (.I(_4100_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9085__A1 (.I(_1382_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9085__A2 (.I(_4113_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9086__A1 (.I(_4041_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9086__B (.I(\as2650.psl[1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9087__C (.I(_3249_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9088__A1 (.I(_1523_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9088__A2 (.I(_0339_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9088__A3 (.I(_4062_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9089__A1 (.I(_1319_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9089__A2 (.I(_2925_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9090__A1 (.I(_4065_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9091__I (.I(_4121_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9092__A1 (.I(_1706_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9092__A2 (.I(_4028_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9093__A1 (.I(_0944_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9093__A2 (.I(_4113_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9094__A1 (.I(_1588_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9094__A2 (.I(_4113_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9095__B (.I(net27));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9096__C (.I(_3249_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9097__A1 (.I(_2373_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9097__A2 (.I(_3144_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9097__B (.I(_4121_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9098__A1 (.I(\as2650.psu[4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9100__A2 (.I(_4129_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9101__B (.I(_3619_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9102__A1 (.I(_3132_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9102__A2 (.I(_4121_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9103__A1 (.I(\as2650.psu[3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9104__A1 (.I(_3133_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9104__A2 (.I(_4028_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9106__B (.I(_1302_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9108__CLK (.I(clknet_leaf_68_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9109__CLK (.I(clknet_leaf_68_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9110__CLK (.I(clknet_leaf_68_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9111__CLK (.I(clknet_leaf_68_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9112__CLK (.I(clknet_leaf_68_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9113__CLK (.I(clknet_leaf_67_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9114__CLK (.I(clknet_leaf_67_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9115__CLK (.I(clknet_leaf_38_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9117__CLK (.I(clknet_leaf_41_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9118__CLK (.I(clknet_leaf_39_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9119__CLK (.I(clknet_leaf_38_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9120__CLK (.I(clknet_leaf_38_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9121__CLK (.I(clknet_leaf_39_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9123__CLK (.I(clknet_leaf_58_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9126__CLK (.I(clknet_leaf_59_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9127__CLK (.I(clknet_leaf_58_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9128__CLK (.I(clknet_leaf_58_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9129__CLK (.I(clknet_leaf_58_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9130__CLK (.I(clknet_leaf_58_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9131__CLK (.I(clknet_leaf_49_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9132__CLK (.I(clknet_leaf_56_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9134__CLK (.I(clknet_leaf_56_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9135__CLK (.I(clknet_leaf_58_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9136__CLK (.I(clknet_leaf_58_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9137__CLK (.I(clknet_leaf_46_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9138__CLK (.I(clknet_leaf_46_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9139__CLK (.I(clknet_leaf_46_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9140__CLK (.I(clknet_leaf_46_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9141__CLK (.I(clknet_leaf_67_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9142__CLK (.I(clknet_leaf_67_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9143__CLK (.I(clknet_leaf_67_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9146__CLK (.I(clknet_leaf_15_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9147__CLK (.I(clknet_leaf_15_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9148__CLK (.I(clknet_leaf_15_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9149__CLK (.I(clknet_leaf_15_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9150__CLK (.I(clknet_leaf_15_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9151__CLK (.I(clknet_leaf_15_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9152__CLK (.I(clknet_leaf_16_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9153__CLK (.I(clknet_leaf_16_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9156__CLK (.I(clknet_leaf_56_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9158__CLK (.I(clknet_leaf_56_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9159__CLK (.I(clknet_leaf_58_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9160__CLK (.I(clknet_leaf_58_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9161__CLK (.I(clknet_3_4_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9162__CLK (.I(clknet_leaf_45_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9162__D (.I(_0055_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9163__CLK (.I(clknet_leaf_48_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9164__CLK (.I(clknet_leaf_48_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9165__CLK (.I(clknet_leaf_48_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9166__CLK (.I(clknet_leaf_48_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9167__CLK (.I(clknet_leaf_49_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9168__CLK (.I(clknet_leaf_48_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9169__CLK (.I(clknet_leaf_48_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9170__CLK (.I(clknet_leaf_60_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9171__CLK (.I(clknet_leaf_60_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9172__CLK (.I(clknet_leaf_60_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9173__CLK (.I(clknet_leaf_60_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9174__CLK (.I(clknet_leaf_60_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9175__CLK (.I(clknet_leaf_60_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9176__CLK (.I(clknet_leaf_59_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9177__D (.I(_0070_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9178__CLK (.I(clknet_leaf_73_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9178__D (.I(_0071_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9179__CLK (.I(clknet_leaf_9_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9183__CLK (.I(clknet_leaf_74_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9184__CLK (.I(clknet_leaf_69_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9185__CLK (.I(clknet_leaf_73_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9186__CLK (.I(clknet_leaf_73_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9187__CLK (.I(clknet_leaf_65_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9188__CLK (.I(clknet_leaf_69_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9189__CLK (.I(clknet_leaf_65_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9190__CLK (.I(clknet_leaf_65_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9191__CLK (.I(clknet_leaf_47_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9192__CLK (.I(clknet_leaf_48_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9193__CLK (.I(clknet_leaf_48_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9194__CLK (.I(clknet_leaf_48_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9195__CLK (.I(clknet_leaf_47_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9196__CLK (.I(clknet_leaf_47_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9197__CLK (.I(clknet_leaf_47_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9198__CLK (.I(clknet_leaf_46_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9199__CLK (.I(clknet_leaf_47_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9200__CLK (.I(clknet_leaf_60_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9201__CLK (.I(clknet_leaf_60_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9202__CLK (.I(clknet_leaf_47_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9203__CLK (.I(clknet_leaf_47_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9204__CLK (.I(clknet_leaf_46_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9205__CLK (.I(clknet_leaf_74_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9206__CLK (.I(clknet_leaf_73_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9207__CLK (.I(clknet_leaf_77_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9208__CLK (.I(clknet_leaf_77_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9210__CLK (.I(clknet_leaf_77_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9211__CLK (.I(clknet_leaf_76_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9213__CLK (.I(clknet_leaf_56_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9214__CLK (.I(clknet_leaf_41_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9215__CLK (.I(clknet_leaf_41_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9216__CLK (.I(clknet_leaf_41_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9218__CLK (.I(clknet_leaf_56_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9219__CLK (.I(clknet_leaf_54_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9220__CLK (.I(clknet_leaf_40_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9221__CLK (.I(clknet_leaf_37_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9222__CLK (.I(clknet_leaf_40_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9223__CLK (.I(clknet_leaf_40_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9224__CLK (.I(clknet_leaf_39_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9225__CLK (.I(clknet_leaf_55_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9226__CLK (.I(clknet_leaf_37_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9228__CLK (.I(clknet_leaf_40_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9229__CLK (.I(clknet_leaf_62_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9232__CLK (.I(clknet_leaf_63_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9233__CLK (.I(clknet_3_0_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9234__CLK (.I(clknet_leaf_62_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9235__CLK (.I(clknet_leaf_62_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9237__CLK (.I(clknet_leaf_55_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9238__CLK (.I(clknet_leaf_39_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9239__CLK (.I(clknet_leaf_39_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9240__CLK (.I(clknet_leaf_38_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9241__CLK (.I(clknet_leaf_55_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9242__CLK (.I(clknet_leaf_55_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9243__CLK (.I(clknet_leaf_55_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9244__CLK (.I(clknet_leaf_39_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9245__CLK (.I(clknet_3_0_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9246__CLK (.I(clknet_leaf_62_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9247__CLK (.I(clknet_leaf_62_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9248__CLK (.I(clknet_leaf_63_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9249__CLK (.I(clknet_3_1_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9251__CLK (.I(clknet_leaf_63_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9252__CLK (.I(clknet_leaf_63_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9253__CLK (.I(clknet_leaf_55_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9254__CLK (.I(clknet_leaf_50_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9255__CLK (.I(clknet_leaf_50_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9256__CLK (.I(clknet_leaf_44_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9257__CLK (.I(clknet_leaf_55_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9258__CLK (.I(clknet_leaf_56_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9259__CLK (.I(clknet_leaf_55_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9260__CLK (.I(clknet_leaf_50_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9261__CLK (.I(clknet_leaf_54_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9262__CLK (.I(clknet_leaf_51_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9263__CLK (.I(clknet_leaf_52_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9264__CLK (.I(clknet_leaf_52_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9265__CLK (.I(clknet_leaf_54_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9266__CLK (.I(clknet_leaf_54_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9267__CLK (.I(clknet_leaf_54_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9268__CLK (.I(clknet_leaf_52_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9270__CLK (.I(clknet_leaf_12_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9272__CLK (.I(clknet_leaf_12_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9273__CLK (.I(clknet_leaf_12_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9276__CLK (.I(clknet_3_2_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9279__CLK (.I(clknet_3_3_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9279__D (.I(_0172_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9280__CLK (.I(clknet_leaf_26_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9281__CLK (.I(clknet_leaf_26_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9281__D (.I(_0174_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9282__CLK (.I(clknet_leaf_26_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9283__CLK (.I(clknet_leaf_26_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9284__CLK (.I(clknet_leaf_26_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9285__CLK (.I(clknet_leaf_27_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9286__CLK (.I(clknet_leaf_27_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9287__CLK (.I(clknet_leaf_27_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9288__CLK (.I(clknet_leaf_27_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9291__CLK (.I(clknet_leaf_31_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9292__CLK (.I(clknet_leaf_31_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9294__CLK (.I(clknet_leaf_25_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9297__CLK (.I(clknet_leaf_3_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9299__CLK (.I(clknet_leaf_1_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9300__CLK (.I(clknet_leaf_1_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9301__CLK (.I(clknet_leaf_1_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9302__CLK (.I(clknet_leaf_1_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9304__CLK (.I(clknet_3_0_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9305__CLK (.I(clknet_3_3_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9308__CLK (.I(clknet_leaf_18_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9309__CLK (.I(clknet_leaf_16_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9310__CLK (.I(clknet_leaf_18_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9311__CLK (.I(clknet_3_3_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9312__CLK (.I(clknet_leaf_18_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9313__CLK (.I(clknet_leaf_18_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9314__CLK (.I(clknet_leaf_9_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9315__CLK (.I(clknet_leaf_24_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9315__D (.I(_0208_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9316__CLK (.I(clknet_3_2_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9316__D (.I(_0209_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9317__CLK (.I(clknet_leaf_25_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9318__CLK (.I(clknet_leaf_30_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9318__D (.I(_0211_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9319__CLK (.I(clknet_3_6_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9319__D (.I(_0212_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9320__CLK (.I(clknet_leaf_31_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9320__D (.I(_0213_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9321__CLK (.I(clknet_leaf_31_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9321__D (.I(_0214_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9323__CLK (.I(clknet_leaf_24_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9325__CLK (.I(clknet_leaf_30_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9326__CLK (.I(clknet_3_6_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9327__CLK (.I(clknet_3_7_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9328__CLK (.I(clknet_3_7_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9328__D (.I(_0221_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9329__CLK (.I(clknet_3_6_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9330__CLK (.I(clknet_leaf_80_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9330__D (.I(_0223_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9331__CLK (.I(clknet_leaf_80_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9331__D (.I(_0224_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9332__CLK (.I(clknet_leaf_80_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9332__D (.I(_0225_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9333__CLK (.I(clknet_leaf_80_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9333__D (.I(_0226_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9334__CLK (.I(clknet_leaf_80_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9334__D (.I(_0227_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9335__CLK (.I(clknet_leaf_80_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9335__D (.I(_0228_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9336__CLK (.I(clknet_3_0_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9336__D (.I(_0229_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9337__CLK (.I(clknet_leaf_77_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9337__D (.I(_0230_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9338__CLK (.I(clknet_leaf_39_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9339__CLK (.I(clknet_leaf_51_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9340__CLK (.I(clknet_leaf_50_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9341__CLK (.I(clknet_leaf_51_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9342__CLK (.I(clknet_leaf_38_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9343__CLK (.I(clknet_leaf_38_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9344__CLK (.I(clknet_leaf_37_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9345__CLK (.I(clknet_leaf_52_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9346__CLK (.I(clknet_leaf_37_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9347__CLK (.I(clknet_leaf_40_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9348__CLK (.I(clknet_leaf_41_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9349__CLK (.I(clknet_leaf_51_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9351__CLK (.I(clknet_leaf_38_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9352__CLK (.I(clknet_leaf_38_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9353__CLK (.I(clknet_leaf_44_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9354__CLK (.I(clknet_leaf_59_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9355__CLK (.I(clknet_leaf_60_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9356__CLK (.I(clknet_leaf_59_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9357__CLK (.I(clknet_leaf_60_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9358__CLK (.I(clknet_leaf_59_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9359__CLK (.I(clknet_leaf_59_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9360__CLK (.I(clknet_leaf_59_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9361__CLK (.I(clknet_leaf_74_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9362__CLK (.I(clknet_leaf_69_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9363__CLK (.I(clknet_leaf_69_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9364__CLK (.I(clknet_leaf_73_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9365__CLK (.I(clknet_3_4_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9366__CLK (.I(clknet_leaf_68_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9367__CLK (.I(clknet_leaf_68_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9368__CLK (.I(clknet_leaf_65_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9369__CLK (.I(clknet_leaf_74_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9370__CLK (.I(clknet_leaf_76_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9371__CLK (.I(clknet_leaf_76_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9372__CLK (.I(clknet_leaf_76_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9373__CLK (.I(clknet_leaf_74_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9374__CLK (.I(clknet_leaf_77_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9376__CLK (.I(clknet_leaf_74_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9377__CLK (.I(clknet_leaf_9_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9379__CLK (.I(clknet_leaf_45_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9379__D (.I(_0272_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9380__CLK (.I(clknet_leaf_44_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9380__D (.I(_0273_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9381__CLK (.I(clknet_leaf_44_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9381__D (.I(_0274_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9382__CLK (.I(clknet_3_2_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9383__CLK (.I(clknet_leaf_3_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9384__CLK (.I(clknet_leaf_3_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9384__D (.I(_0277_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9385__D (.I(_0278_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9386__CLK (.I(clknet_leaf_3_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9386__D (.I(_0279_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__9388__CLK (.I(clknet_3_1_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_0_wb_clk_i_I (.I(wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_3_0_0_wb_clk_i_I (.I(clknet_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_3_1_0_wb_clk_i_I (.I(clknet_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_3_2_0_wb_clk_i_I (.I(clknet_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_3_3_0_wb_clk_i_I (.I(clknet_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_3_4_0_wb_clk_i_I (.I(clknet_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_3_5_0_wb_clk_i_I (.I(clknet_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_3_6_0_wb_clk_i_I (.I(clknet_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_3_7_0_wb_clk_i_I (.I(clknet_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_11_wb_clk_i_I (.I(clknet_3_2_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_12_wb_clk_i_I (.I(clknet_3_2_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_14_wb_clk_i_I (.I(clknet_3_2_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_15_wb_clk_i_I (.I(clknet_3_2_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_16_wb_clk_i_I (.I(clknet_3_3_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_18_wb_clk_i_I (.I(clknet_3_3_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_1_wb_clk_i_I (.I(clknet_3_0_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_20_wb_clk_i_I (.I(clknet_3_3_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_23_wb_clk_i_I (.I(clknet_3_3_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_24_wb_clk_i_I (.I(clknet_3_6_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_25_wb_clk_i_I (.I(clknet_3_6_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_26_wb_clk_i_I (.I(clknet_opt_1_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_27_wb_clk_i_I (.I(clknet_3_6_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_28_wb_clk_i_I (.I(clknet_3_6_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_29_wb_clk_i_I (.I(clknet_3_6_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_2_wb_clk_i_I (.I(clknet_3_0_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_30_wb_clk_i_I (.I(clknet_3_6_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_31_wb_clk_i_I (.I(clknet_3_6_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_36_wb_clk_i_I (.I(clknet_3_7_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_37_wb_clk_i_I (.I(clknet_3_7_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_38_wb_clk_i_I (.I(clknet_3_7_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_39_wb_clk_i_I (.I(clknet_3_7_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_3_wb_clk_i_I (.I(clknet_3_2_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_40_wb_clk_i_I (.I(clknet_3_7_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_41_wb_clk_i_I (.I(clknet_3_7_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_42_wb_clk_i_I (.I(clknet_3_7_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_44_wb_clk_i_I (.I(clknet_3_5_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_45_wb_clk_i_I (.I(clknet_3_5_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_46_wb_clk_i_I (.I(clknet_3_4_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_47_wb_clk_i_I (.I(clknet_3_5_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_48_wb_clk_i_I (.I(clknet_3_5_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_49_wb_clk_i_I (.I(clknet_3_5_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_50_wb_clk_i_I (.I(clknet_3_5_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_51_wb_clk_i_I (.I(clknet_3_7_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_52_wb_clk_i_I (.I(clknet_3_5_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_53_wb_clk_i_I (.I(clknet_3_5_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_54_wb_clk_i_I (.I(clknet_3_5_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_55_wb_clk_i_I (.I(clknet_3_5_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_56_wb_clk_i_I (.I(clknet_3_5_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_57_wb_clk_i_I (.I(clknet_3_5_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_58_wb_clk_i_I (.I(clknet_3_5_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_59_wb_clk_i_I (.I(clknet_3_5_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_5_wb_clk_i_I (.I(clknet_3_1_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_60_wb_clk_i_I (.I(clknet_3_5_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_61_wb_clk_i_I (.I(clknet_3_5_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_62_wb_clk_i_I (.I(clknet_3_4_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_63_wb_clk_i_I (.I(clknet_3_4_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_64_wb_clk_i_I (.I(clknet_3_4_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_65_wb_clk_i_I (.I(clknet_3_4_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_66_wb_clk_i_I (.I(clknet_3_4_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_67_wb_clk_i_I (.I(clknet_3_4_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_68_wb_clk_i_I (.I(clknet_3_4_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_69_wb_clk_i_I (.I(clknet_3_4_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_6_wb_clk_i_I (.I(clknet_3_1_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_71_wb_clk_i_I (.I(clknet_3_4_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_73_wb_clk_i_I (.I(clknet_3_1_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_74_wb_clk_i_I (.I(clknet_3_1_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_75_wb_clk_i_I (.I(clknet_3_1_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_76_wb_clk_i_I (.I(clknet_3_1_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_77_wb_clk_i_I (.I(clknet_3_1_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_80_wb_clk_i_I (.I(clknet_3_0_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_8_wb_clk_i_I (.I(clknet_3_3_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_9_wb_clk_i_I (.I(clknet_3_3_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_opt_1_0_wb_clk_i_I (.I(clknet_3_6_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout51_I (.I(net25));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout52_I (.I(net40));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout53_I (.I(net38));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout54_I (.I(net35));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input10_I (.I(io_in[9]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input1_I (.I(io_in[10]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input2_I (.I(io_in[11]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input3_I (.I(io_in[12]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input4_I (.I(io_in[13]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input5_I (.I(io_in[33]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input6_I (.I(io_in[5]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input7_I (.I(io_in[6]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input8_I (.I(io_in[7]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input9_I (.I(io_in[8]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output14_I (.I(net14));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output15_I (.I(net15));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output16_I (.I(net16));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output17_I (.I(net17));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output18_I (.I(net18));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output21_I (.I(net21));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output23_I (.I(net23));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output24_I (.I(net24));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output25_I (.I(net25));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output26_I (.I(net26));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output27_I (.I(net27));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output31_I (.I(net31));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output33_I (.I(net33));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output34_I (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output35_I (.I(net35));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output36_I (.I(net36));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output37_I (.I(net37));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output38_I (.I(net38));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output39_I (.I(net39));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output40_I (.I(net40));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1014 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_1025 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1029 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_1037 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_1045 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1049 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1066 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1073 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_1077 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_1094 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_1110 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1118 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1154 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_1183 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1187 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1189 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_1208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1222 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1224 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1227 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1257 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1259 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1262 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1264 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1294 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_1297 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1329 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_1332 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1364 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_1367 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1391 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1398 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_1402 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1434 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_1437 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1469 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_1472 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1504 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_1507 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1539 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_1542 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1574 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_1577 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_569 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_585 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_593 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_629 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_664 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_699 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_734 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_769 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_788 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_792 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_799 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_803 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_839 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_874 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_884 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_892 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_908 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_944 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_979 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_982 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_100_10 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_100_1018 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_1026 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_103 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_100_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_1037 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_1045 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_1057 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_1068 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_1072 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_100_1076 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_100_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_100_1092 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_100_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_1106 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_1110 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_100_1114 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_1118 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_100_1125 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_114 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_100_1141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_1149 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_100_1156 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_100_1164 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_1168 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_1179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_1183 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_1187 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_1191 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_1198 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_1204 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_1210 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_100_1214 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_1224 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_1228 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_100_1232 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_1236 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_1238 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_100_1274 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_1282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_1293 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_100_1309 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_100_1318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_132 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_1328 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_1334 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_100_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_100_1380 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_1389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_100_1393 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_14 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_100_1406 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_143 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_100_1438 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_100_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_100_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_100_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_155 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_100_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_100_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_161 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_100_195 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_100_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_204 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_211 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_222 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_23 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_100_253 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_263 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_27 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_271 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_100_275 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_287 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_291 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_297 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_305 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_100_31 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_313 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_100_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_100_337 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_347 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_351 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_359 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_367 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_100_371 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_398 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_100_40 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_100_402 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_100_434 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_44 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_100_450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_458 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_100_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_100_47 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_477 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_100_481 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_497 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_100_501 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_51 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_100_517 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_100_525 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_529 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_100_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_55 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_59 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_100_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_100_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_100_621 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_100_629 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_63 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_633 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_100_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_67 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_100_670 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_100_679 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_743 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_100_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_755 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_757 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_764 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_100_768 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_77 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_100_800 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_100_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_850 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_853 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_865 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_869 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_873 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_100_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_885 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_100_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_100_921 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_93 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_937 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_941 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_100_949 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_100_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_100_968 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_972 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_975 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_982 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_100_986 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_1014 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_101_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_1032 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_1034 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_1037 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_1041 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_1045 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_101_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_1057 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_101_1061 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_1074 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_1076 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_101_1083 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_1091 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_1094 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_1098 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_101_1108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_111 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_101_1118 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_1124 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_101_1127 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_1142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_101_1150 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_101_1158 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_1162 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_1178 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_1190 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_1194 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_1196 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_1212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_1216 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_101_1220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_1230 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_1242 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_1246 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_101_1250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_1254 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_1261 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_101_1265 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_101_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_101_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_1290 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_1298 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_101_1302 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_101_1318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_101_1326 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_1330 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_1334 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_1357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_101_1361 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_1393 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_101_1397 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_140 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_101_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_101_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_101_147 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_101_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_101_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_153 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_101_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_101_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_101_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_184 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_191 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_197 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_101_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_204 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_101_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_22 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_221 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_101_225 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_229 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_238 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_101_242 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_101_25 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_101_258 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_262 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_101_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_310 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_101_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_328 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_33 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_332 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_336 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_101_340 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_101_348 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_36 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_364 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_368 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_101_372 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_101_388 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_394 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_399 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_101_403 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_101_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_423 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_101_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_43 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_101_434 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_101_466 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_101_482 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_488 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_101_491 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_495 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_101_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_51 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_101_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_101_547 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_101_55 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_101_553 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_101_561 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_101_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_586 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_59 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_593 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_101_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_101_613 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_62 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_101_621 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_625 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_627 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_636 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_101_644 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_101_660 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_666 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_674 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_685 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_101_689 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_101_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_101_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_76 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_101_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_785 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_792 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_101_796 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_101_812 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_101_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_101_824 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_101_840 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_848 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_866 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_878 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_101_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_101_902 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_910 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_101_928 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_93 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_101_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_976 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_980 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_101_984 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_992 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_101_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_102_1006 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_1014 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_1020 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_1035 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_1047 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_102_1055 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_1071 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_102_1077 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_1093 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_1097 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_1106 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_1113 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_1117 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_112 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_1121 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_1125 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_1137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_114 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_1141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_1144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_102_1152 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_117 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_1182 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_1186 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_1193 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_1197 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_1204 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_1216 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_1220 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_1224 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_1228 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_124 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_1240 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_1247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_1251 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_102_1255 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_102_1287 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_1303 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_1305 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_102_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_1331 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_1335 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_1349 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_1357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_1361 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_1365 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_1369 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_1373 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_102_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_1394 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_1398 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_1400 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_1403 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_1413 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_1426 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_1428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_1437 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_102_1441 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_1449 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_1453 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_102_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_102_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_155 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_102_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_163 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_167 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_169 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_186 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_192 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_102_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_202 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_102_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_216 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_224 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_228 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_102_232 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_102_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_290 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_102_298 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_334 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_342 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_102_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_358 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_362 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_364 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_370 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_374 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_102_378 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_386 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_394 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_400 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_404 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_102_408 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_420 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_430 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_438 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_102_442 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_458 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_469 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_495 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_102_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_507 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_537 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_541 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_551 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_565 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_571 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_575 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_579 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_581 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_584 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_591 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_102_595 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_60 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_102_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_613 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_102_616 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_102_648 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_102_664 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_672 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_102_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_68 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_102_708 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_716 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_720 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_722 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_729 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_102_733 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_741 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_102_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_102_763 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_773 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_78 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_784 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_790 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_794 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_814 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_821 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_825 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_102_832 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_866 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_102_870 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_102_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_905 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_909 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_923 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_933 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_937 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_941 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_102_945 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_97 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_972 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_976 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_986 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_102_990 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_103_1004 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_103_1014 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_103_103 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_103_1030 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_1038 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_1040 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_1043 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_1047 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_1051 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_103_1059 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_1063 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_103_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_103_1075 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_1079 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_1109 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_1113 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_103_1117 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_1125 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_103_1129 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_1133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_103_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_1144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_1152 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_1154 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_103_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_1163 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_1171 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_1180 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_1184 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_103_1188 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_103_119 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_1195 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_103_1199 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_103_1212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_1228 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_123 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_1232 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_1240 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_1242 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_103_1245 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_126 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_103_1261 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_103_1269 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_1276 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_103_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_103_1286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_1292 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_1299 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_103_1303 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_1307 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_132 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_1337 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_1341 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_103_1345 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_103_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_1367 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_103_1374 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_103_1382 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_1389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_1393 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_103_1403 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_103_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_1438 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_1440 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_103_1443 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_1451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_103_1460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_103_1476 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_103_1484 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_1488 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_103_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_103_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_103_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_103_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_195 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_103_199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_103_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_203 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_224 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_231 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_103_235 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_254 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_258 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_103_26 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_260 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_263 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_270 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_103_274 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_103_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_30 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_32 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_328 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_342 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_35 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_353 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_103_364 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_368 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_103_375 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_39 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_103_391 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_399 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_401 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_404 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_411 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_103_415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_423 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_103_432 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_103_47 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_103_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_103_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_103_547 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_103_553 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_103_561 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_565 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_57 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_103_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_578 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_581 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_103_585 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_59 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_103_601 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_607 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_614 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_62 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_624 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_103_628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_636 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_103_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_103_649 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_655 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_665 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_103_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_103_701 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_103_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_103_728 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_103_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_738 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_103_751 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_103_767 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_103_775 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_779 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_785 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_788 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_79 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_103_792 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_103_826 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_103_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_850 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_103_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_103_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_103_928 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_94 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_96 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_962 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_968 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_972 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_976 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_103_980 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_103_988 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_99 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_992 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_103_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_100 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_1008 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_1011 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_1020 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_104_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_104_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_1047 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_1056 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_1065 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_1069 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_104_1073 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_104_1089 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_1097 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_104_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_1110 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_1113 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_1125 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_1129 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_104_1133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_1137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_1144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_104_115 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_1155 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_1159 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_1163 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_104_1167 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_1184 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_1188 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_104_1196 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_104_1212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_104_1220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_1224 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_1228 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_123 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_1232 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_104_1251 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_1259 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_1262 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_104_1274 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_1286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_1296 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_104_1300 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_104_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_1331 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_1339 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_1350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_1354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_104_1358 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_1362 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_1366 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_104_1389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_1397 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_1399 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_104_1402 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_104_1418 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_104_1426 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_1430 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_1432 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_1435 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_104_1439 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_1463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_104_1467 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_104_1499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_104_1515 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_1523 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_104_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_104_154 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_104_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_104_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_164 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_104_182 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_192 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_104_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_200 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_104_204 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_214 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_104_217 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_233 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_237 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_104_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_261 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_269 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_271 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_274 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_290 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_294 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_296 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_104_303 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_307 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_310 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_323 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_326 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_337 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_341 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_104_345 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_104_361 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_365 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_104_369 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_104_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_104_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_104_408 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_104_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_420 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_423 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_104_431 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_445 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_449 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_104_453 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_471 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_104_475 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_104_507 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_515 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_104_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_104_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_550 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_552 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_579 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_589 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_104_593 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_599 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_61 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_104_624 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_630 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_104_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_65 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_67 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_104_670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_104_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_104_684 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_690 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_694 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_104_710 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_742 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_104_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_104_779 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_104_787 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_79 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_791 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_104_794 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_104_810 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_814 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_104_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_87 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_104_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_104_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_91 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_93 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_104_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_104_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_104_992 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_1004 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_1008 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_105_102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_105_1020 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_105_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_1034 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_1038 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_1050 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_1054 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_1063 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_105_1070 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_105_1078 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_1084 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_1088 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_1100 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_1104 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_105_1108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_105_1116 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_1120 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_1128 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_105_1132 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_1141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_1143 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_105_1149 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_1161 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_1165 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_1167 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_105_118 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_1182 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_1186 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_1190 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_1194 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_1196 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_1205 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_105_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_1225 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_1227 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_1230 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_1234 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_1250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_1254 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_1258 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_126 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_105_1262 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_128 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_105_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_1284 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_1288 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_105_1292 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_131 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_105_1324 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_1330 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_105_1345 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_105_1359 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_105_1369 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_105_1385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_1391 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_1401 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_1405 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_1409 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_1413 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_1417 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_105_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_105_1430 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_1436 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_105_1444 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_147 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_105_1476 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_105_1484 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_1488 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_105_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_151 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_153 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_105_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_156 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_105_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_160 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_105_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_105_191 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_105_197 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_105_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_105_223 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_231 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_105_235 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_105_256 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_105_26 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_260 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_262 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_268 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_105_272 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_105_280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_105_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_302 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_105_305 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_313 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_32 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_328 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_105_336 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_363 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_105_367 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_38 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_105_383 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_391 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_394 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_398 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_410 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_105_414 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_105_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_105_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_105_444 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_448 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_458 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_105_462 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_494 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_105_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_105_505 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_509 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_512 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_516 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_529 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_105_533 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_566 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_574 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_584 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_105_63 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_636 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_105_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_649 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_653 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_663 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_105_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_67 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_105_683 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_693 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_105_715 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_105_731 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_739 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_105_743 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_775 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_777 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_105_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_105_792 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_798 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_105_808 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_81 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_816 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_819 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_823 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_838 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_105_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_850 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_105_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_870 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_873 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_883 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_887 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_105_891 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_105_909 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_105_917 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_921 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_105_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_105_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_961 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_965 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_969 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_981 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_985 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_105_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_105_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_106_1002 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_1011 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_106_1015 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_106_1023 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_1027 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_106_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_106_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_1043 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_1047 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_1059 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_1063 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_106_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_1071 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_1074 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_1082 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_106_1090 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_1098 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_106_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_106_111 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_106_1110 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_1114 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_1124 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_1128 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_1137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_1141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_1143 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_1146 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_1150 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_1154 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_1158 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_1162 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_106_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_106_1176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_106_1184 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_1188 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_1190 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_1193 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_106_1197 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_106_1229 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_106_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_106_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_106_1260 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_106_127 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_1270 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_106_1278 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_1310 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_106_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_106_1331 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_1335 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_1337 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_106_1352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_1356 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_1358 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_1361 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_106_1365 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_1381 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_1389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_140 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_1402 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_1412 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_1420 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_106_1424 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_1440 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_1444 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_1446 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_1453 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_106_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_147 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_106_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_106_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_106_154 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_106_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_106_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_164 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_186 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_106_193 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_106_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_202 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_106_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_106_214 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_218 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_221 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_106_233 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_239 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_106_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_106_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_268 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_106_284 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_106_292 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_296 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_298 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_106_304 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_106_312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_316 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_323 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_326 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_106_330 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_358 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_360 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_366 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_106_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_370 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_106_374 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_106_382 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_386 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_399 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_406 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_106_410 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_106_442 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_450 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_106_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_458 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_106_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_467 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_469 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_106_47 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_472 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_476 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_478 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_106_481 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_106_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_106_503 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_509 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_106_513 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_529 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_106_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_55 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_106_550 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_554 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_556 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_59 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_593 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_601 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_63 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_106_635 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_651 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_654 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_658 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_665 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_67 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_672 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_106_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_106_708 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_106_716 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_720 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_722 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_725 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_729 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_106_741 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_106_750 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_106_758 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_106_764 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_106_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_788 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_79 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_796 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_106_800 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_106_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_834 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_838 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_106_857 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_106_873 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_106_881 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_885 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_106_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_897 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_901 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_106_905 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_106_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_930 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_933 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_106_941 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_106_949 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_106_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_970 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_106_978 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_106_994 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_1012 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_1014 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_107_1020 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_107_1030 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_107_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_1062 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_1073 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_1077 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_1081 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_1085 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_1089 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_1097 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_107_1101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_1105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_1108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_1112 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_1125 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_107_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_1148 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_1156 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_1160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_1162 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_1177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_1181 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_107_1185 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_107_1201 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_1205 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_107_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_1217 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_1220 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_107_1224 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_107_1240 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_1254 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_1258 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_1262 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_107_1270 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_1274 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_107_1287 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_107_1303 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_1311 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_1318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_1324 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_107_1328 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_107_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_107_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_1367 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_1375 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_107_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_1385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_1388 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_107_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_107_1430 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_1436 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_107_1440 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_1455 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_1459 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_107_1463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_107_1479 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_148 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_107_1487 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_107_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_152 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_107_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_156 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_107_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_107_164 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_168 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_107_178 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_184 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_107_188 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_192 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_195 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_107_199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_107_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_107_207 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_211 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_107_227 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_233 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_107_237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_259 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_263 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_267 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_271 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_278 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_107_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_107_294 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_298 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_301 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_313 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_320 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_107_324 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_107_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_107_340 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_107_348 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_107_364 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_396 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_398 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_107_401 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_107_417 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_107_42 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_107_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_107_436 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_440 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_46 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_468 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_107_477 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_483 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_487 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_502 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_506 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_510 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_107_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_53 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_107_537 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_550 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_107_554 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_107_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_566 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_107_57 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_107_584 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_107_616 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_630 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_637 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_107_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_107_649 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_107_65 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_653 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_655 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_107_658 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_107_690 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_107_706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_107_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_107_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_748 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_762 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_77 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_107_770 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_778 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_107_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_787 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_107_790 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_81 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_107_822 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_107_838 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_107_846 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_85 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_850 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_107_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_107_870 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_107_878 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_884 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_887 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_107_89 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_891 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_107_903 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_107_919 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_107_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_93 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_107_961 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_969 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_107_972 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_107_988 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_992 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_107_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_1003 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_108_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_1010 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_108_1014 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_1018 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_1021 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_1038 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_1045 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_108_1049 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_108_1057 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_1061 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_1063 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_108_1066 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_108_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_1082 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_1084 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_108_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_1156 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_1169 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_1179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_1183 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_1187 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_1191 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_108_1195 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_108_1203 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_1207 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_1212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_1220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_1233 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_108_124 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_1246 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_1255 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_1259 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_108_1263 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_128 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_1281 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_1285 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_108_1289 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_1295 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_1299 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_1317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_1329 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_1333 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_1337 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_1341 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_108_1345 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_1349 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_108_1352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_1360 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_108_1363 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_1367 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_1369 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_1372 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_108_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_108_1404 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_1420 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_108_1424 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_108_1432 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_108_1438 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_145 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_108_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_108_1465 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_108_1471 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_108_149 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_108_1503 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_108_1519 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_1523 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_108_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_153 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_108_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_108_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_168 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_182 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_192 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_108_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_108_203 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_108_219 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_108_229 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_245 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_252 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_255 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_259 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_267 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_269 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_272 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_292 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_108_296 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_108_304 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_310 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_328 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_336 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_108_340 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_108_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_108_372 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_388 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_108_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_108_400 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_410 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_108_414 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_108_446 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_452 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_108_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_470 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_474 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_476 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_479 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_108_483 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_487 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_108_500 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_108_516 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_108_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_528 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_536 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_108_543 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_108_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_571 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_575 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_108_579 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_587 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_589 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_108_596 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_600 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_108_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_108_621 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_625 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_628 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_108_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_640 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_642 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_645 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_108_653 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_108_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_108_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_108_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_108_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_108_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_108_755 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_759 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_761 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_108_764 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_108_796 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_108_812 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_108_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_834 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_836 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_839 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_108_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_108_855 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_87 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_108_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_108_905 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_911 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_929 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_108_933 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_108_949 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_962 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_97 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_974 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_978 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_108_982 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_986 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_109_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_109_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_109_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_1058 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_1062 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_109_1078 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_109_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_109_1094 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_1098 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_1100 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_109_1103 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_1119 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_1121 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_1124 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_1144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_1148 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_1152 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_1156 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_109_1160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_1172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_1180 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_1184 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_1188 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_1196 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_109_1200 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_1219 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_109_1227 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_1235 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_124 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_1240 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_1248 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_1258 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_126 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_1262 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_1264 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_1271 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_1275 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_1283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_109_1287 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_109_1303 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_1311 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_1314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_1318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_1322 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_109_1326 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_133 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_109_1342 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_1361 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_1369 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_1373 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_109_1377 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_1390 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_1394 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_1398 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_140 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_109_1402 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_1410 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_1413 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_1417 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_1436 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_109_1444 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_109_1452 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_1456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_146 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_1460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_1464 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_1471 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_109_1482 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_109_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_109_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_109_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_159 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_184 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_188 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_190 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_193 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_109_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_201 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_109_205 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_109_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_109_231 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_235 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_240 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_248 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_109_252 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_109_273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_109_280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_297 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_109_301 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_319 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_109_322 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_109_338 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_109_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_353 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_109_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_109_36 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_109_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_397 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_401 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_411 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_423 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_109_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_109_436 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_442 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_449 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_487 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_491 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_495 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_109_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_515 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_518 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_52 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_522 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_109_526 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_530 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_533 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_109_541 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_109_557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_578 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_593 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_601 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_109_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_61 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_109_613 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_619 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_626 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_109_644 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_65 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_109_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_682 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_109_690 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_109_706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_109_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_109_728 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_109_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_109_736 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_746 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_109_750 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_109_766 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_109_774 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_778 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_109_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_109_81 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_109_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_823 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_830 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_109_834 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_844 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_865 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_109_869 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_109_885 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_891 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_894 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_898 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_908 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_109_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_920 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_109_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_93 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_933 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_935 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_938 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_946 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_948 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_109_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_109_963 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_967 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_969 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_972 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_979 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_109_983 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_991 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_109_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_10_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_10_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_10_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_10_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_10_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_10_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_10_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_10_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_10_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_10_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_10_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_10_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_10_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_10_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_10_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_10_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_10_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_10_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_10_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_10_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_10_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_10_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_10_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_10_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_110_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_1027 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_110_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_110_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_1043 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_1045 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_1048 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_1059 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_1063 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_1065 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_1068 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_110_1072 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_110_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_110_1088 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_110_1096 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_110_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_1106 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_1109 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_1119 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_1123 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_1127 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_1133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_1136 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_1143 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_1153 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_1163 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_110_1167 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_1176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_1180 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_1182 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_1213 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_110_1217 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_110_1233 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_110_124 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_1247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_1259 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_1267 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_1271 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_1275 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_1283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_1296 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_110_1300 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_110_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_110_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_132 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_110_1331 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_1337 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_110_1345 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_110_135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_110_1377 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_1381 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_1389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_1399 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_1409 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_1413 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_110_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_1420 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_110_1424 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_110_1440 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_110_1448 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_1452 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_110_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_110_1465 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_1469 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_110_1473 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_110_150 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_110_1505 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_110_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_110_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_154 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_110_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_157 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_110_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_167 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_175 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_186 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_110_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_200 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_110_204 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_224 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_238 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_245 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_110_253 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_261 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_110_268 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_272 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_110_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_284 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_110_287 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_110_295 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_307 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_110_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_110_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_325 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_110_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_353 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_366 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_110_370 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_110_378 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_382 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_40 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_110_401 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_110_433 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_44 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_110_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_459 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_46 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_110_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_479 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_481 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_49 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_110_490 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_500 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_110_504 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_518 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_530 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_110_537 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_110_553 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_560 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_576 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_110_580 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_584 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_587 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_595 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_110_599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_110_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_110_637 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_64 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_110_653 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_657 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_659 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_662 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_110_670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_110_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_708 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_711 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_721 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_725 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_110_729 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_110_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_755 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_757 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_110_76 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_760 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_767 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_110_771 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_781 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_785 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_799 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_803 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_110_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_110_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_110_850 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_857 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_110_865 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_110_881 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_885 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_110_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_905 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_92 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_94 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_110_963 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_97 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_111_1007 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_1025 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_1029 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_111_1043 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_111_1059 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_1063 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_111_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_111_1083 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_111_1091 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_1097 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_1106 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_1120 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_1124 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_1128 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_1141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_1143 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_111_1154 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_1158 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_116 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_1165 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_111_1175 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_1187 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_1197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_120 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_1201 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_1205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_1225 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_111_1229 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_111_124 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_111_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_1249 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_1253 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_1265 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_1269 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_1283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_1287 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_1289 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_111_1292 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_111_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_1314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_1321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_111_1325 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_1335 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_111_1343 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_1347 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_111_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_1387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_1391 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_1393 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_140 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_1405 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_1417 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_111_1425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_111_1433 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_1437 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_111_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_1441 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_1443 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_1446 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_111_1458 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_111_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_152 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_154 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_111_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_111_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_157 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_161 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_168 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_111_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_184 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_111_188 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_192 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_196 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_111_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_211 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_111_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_111_223 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_227 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_111_231 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_239 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_242 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_111_246 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_111_254 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_111_260 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_264 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_274 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_111_289 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_297 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_299 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_302 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_310 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_111_327 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_111_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_111_343 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_347 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_111_351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_111_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_111_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_111_397 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_401 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_403 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_410 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_111_414 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_111_42 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_111_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_435 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_111_439 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_46 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_111_471 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_475 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_477 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_48 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_494 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_111_502 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_508 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_532 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_111_536 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_545 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_111_549 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_565 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_57 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_111_573 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_577 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_111_584 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_594 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_111_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_618 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_111_622 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_630 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_65 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_656 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_660 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_111_664 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_672 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_674 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_677 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_111_685 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_111_701 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_111_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_111_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_111_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_111_760 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_111_768 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_111_790 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_798 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_802 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_809 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_111_813 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_111_845 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_849 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_111_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_111_862 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_866 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_868 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_111_871 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_887 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_111_890 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_900 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_111_904 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_91 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_920 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_111_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_111_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_973 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_976 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_111_980 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_111_988 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_992 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_999 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_100 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_112_1006 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_1010 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_112_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_1025 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_112_1042 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_112_1058 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_1062 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_1065 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_1073 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_112_1077 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_112_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_1114 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_1126 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_1133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_1137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_1141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_1149 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_1153 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_1155 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_1165 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_1169 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_112_1176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_1180 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_1191 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_1195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_1197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_1208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_1212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_112_1216 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_1232 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_1234 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_1239 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_112_124 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_1256 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_1260 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_1264 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_112_1268 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_112_1276 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_1282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_1290 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_112_1303 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_1311 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_112_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_1319 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_1323 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_1337 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_112_1341 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_112_1361 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_112_1377 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_1381 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_112_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_1390 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_112_1394 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_140 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_1407 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_1411 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_112_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_1437 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_1441 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_112_1460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_112_1468 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_1472 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_1474 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_148 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_1480 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_112_1484 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_150 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_112_1516 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_1524 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_112_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_112_153 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_112_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_112_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_112_169 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_112_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_187 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_112_190 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_198 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_112_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_112_201 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_112_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_213 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_218 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_222 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_229 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_112_233 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_237 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_112_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_257 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_259 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_266 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_112_270 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_112_278 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_112_285 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_293 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_295 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_298 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_112_302 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_112_308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_327 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_112_331 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_112_339 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_343 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_347 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_112_358 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_112_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_112_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_424 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_112_436 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_445 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_112_449 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_112_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_112_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_112_479 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_483 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_485 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_488 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_500 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_112_504 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_508 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_510 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_513 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_517 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_112_53 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_112_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_538 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_112_542 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_550 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_554 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_112_564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_57 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_112_572 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_576 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_112_583 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_592 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_112_599 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_61 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_112_611 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_112_643 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_112_65 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_657 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_112_661 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_671 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_112_679 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_112_711 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_112_727 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_735 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_756 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_112_760 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_112_792 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_112_800 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_804 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_112_81 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_813 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_112_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_85 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_112_850 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_858 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_860 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_863 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_112_867 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_87 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_112_879 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_883 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_112_898 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_902 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_913 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_917 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_112_921 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_96 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_112_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_112_974 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_986 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_112_990 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_100 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_113_1007 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_1011 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_1014 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_1018 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_113_1030 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_113_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_1062 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_1074 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_1082 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_113_1086 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_113_1132 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_1141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_1145 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_1149 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_1153 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_1163 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_1179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_1191 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_1195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_1199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_113_1203 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_113_1212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_113_1220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_1224 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_1231 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_113_1235 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_1245 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_113_1249 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_1257 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_1259 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_113_1262 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_113_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_113_1290 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_113_1306 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_1310 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_1313 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_113_1317 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_113_1333 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_1337 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_1340 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_113_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_1362 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_1366 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_1368 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_1371 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_1375 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_113_1389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_140 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_113_1405 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_113_1413 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_1417 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_113_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_1438 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_1440 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_113_1443 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_1459 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_1462 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_113_1470 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_113_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_113_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_151 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_113_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_113_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_157 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_161 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_186 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_113_196 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_113_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_200 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_113_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_219 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_231 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_238 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_242 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_113_246 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_262 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_113_266 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_274 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_113_293 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_297 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_306 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_113_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_113_337 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_113_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_341 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_113_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_113_373 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_113_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_388 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_395 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_113_399 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_113_415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_423 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_113_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_432 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_440 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_448 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_113_452 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_462 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_113_466 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_113_482 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_113_490 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_494 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_113_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_113_50 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_533 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_540 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_548 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_113_552 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_113_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_578 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_113_58 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_581 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_589 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_591 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_594 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_600 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_603 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_113_615 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_62 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_113_631 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_113_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_651 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_113_658 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_662 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_113_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_113_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_113_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_113_76 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_113_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_113_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_817 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_827 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_113_831 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_84 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_113_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_113_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_86 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_113_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_113_894 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_898 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_113_901 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_917 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_919 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_934 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_938 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_113_942 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_113_958 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_966 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_970 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_979 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_113_983 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_991 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_113_999 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_114_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_103 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_114_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_114_1063 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_1071 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_1073 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_114_1076 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_114_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_1092 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_1114 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_1118 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_114_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_1128 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_1132 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_1136 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_114_1140 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_1148 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_1152 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_1156 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_1160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_1164 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_1168 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_1177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_1181 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_1185 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_1189 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_1191 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_1194 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_1198 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_114_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_114_1210 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_114_1218 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_1222 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_1224 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_114_1227 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_1231 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_1234 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_1257 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_114_1261 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_1279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_1282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_114_1286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_1302 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_1311 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_1328 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_114_1332 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_1350 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_114_1354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_114_1370 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_114_1378 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_1382 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_114_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_1402 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_1406 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_1414 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_1418 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_114_1426 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_114_1442 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_114_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_114_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_114_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_114_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_153 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_114_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_114_157 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_114_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_114_173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_184 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_114_188 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_192 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_195 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_114_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_220 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_114_227 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_233 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_239 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_242 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_114_259 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_269 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_114_277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_281 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_290 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_294 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_301 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_303 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_309 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_316 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_326 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_114_330 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_334 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_336 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_339 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_364 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_114_368 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_114_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_114_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_388 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_403 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_407 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_114_411 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_424 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_432 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_114_436 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_114_442 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_114_45 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_458 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_114_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_114_479 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_487 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_49 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_495 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_114_503 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_51 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_114_519 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_114_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_114_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_538 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_114_542 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_114_558 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_566 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_568 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_114_571 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_58 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_114_587 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_591 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_593 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_600 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_608 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_114_616 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_62 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_114_624 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_631 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_639 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_114_643 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_659 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_114_663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_671 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_114_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_114_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_114_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_114_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_781 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_788 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_114_792 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_114_808 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_114_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_826 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_828 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_831 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_844 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_848 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_852 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_856 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_86 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_114_860 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_114_876 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_884 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_114_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_114_921 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_929 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_933 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_937 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_95 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_114_951 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_955 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_114_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_99 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_1014 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_115_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_115_1040 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_1048 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_1051 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_1059 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_1061 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_115_1074 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_1082 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_1085 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_1089 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_1106 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_1110 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_1114 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_1118 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_115_112 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_1128 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_115_1132 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_1141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_1143 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_115_1146 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_1152 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_1161 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_1165 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_115_1169 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_1185 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_115_1188 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_1195 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_115_1199 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_1203 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_1220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_1224 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_1226 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_115_1235 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_1243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_1249 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_115_1253 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_115_1261 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_1267 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_115_128 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_1283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_1285 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_115_1298 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_115_1306 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_1310 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_115_1314 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_115_1330 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_1336 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_1354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_1358 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_115_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_1360 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_1363 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_115_1373 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_140 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_1407 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_115_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_115_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_1428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_115_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_1442 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_1449 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_115_1453 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_115_1461 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_1467 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_1471 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_1481 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_115_1485 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_1489 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_115_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_115_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_115_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_115_160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_115_178 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_182 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_115_186 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_192 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_115_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_223 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_225 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_228 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_240 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_251 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_115_255 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_115_263 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_267 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_269 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_272 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_293 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_115_297 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_303 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_305 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_322 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_115_330 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_115_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_115_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_366 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_115_370 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_38 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_115_402 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_115_418 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_115_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_436 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_115_444 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_452 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_115_455 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_115_470 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_115_480 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_506 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_510 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_522 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_543 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_115_547 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_551 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_561 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_577 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_579 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_582 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_115_593 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_607 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_115_611 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_62 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_115_627 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_635 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_115_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_653 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_115_657 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_115_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_681 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_684 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_692 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_115_696 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_115_704 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_708 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_725 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_729 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_115_733 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_115_749 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_115_757 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_76 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_768 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_115_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_115_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_115_80 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_115_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_115_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_115_862 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_866 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_868 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_115_871 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_115_903 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_115_911 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_915 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_115_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_115_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_115_941 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_949 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_115_964 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_115_980 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_115_988 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_992 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_115_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_100 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_1005 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_1009 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_1019 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_1026 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_116_1034 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_1038 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_1040 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_1043 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_116_1047 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_116_1079 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_1093 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_1097 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_1105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_116_1113 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_116_1121 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_1125 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_1128 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_1132 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_1144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_1161 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_116_1165 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_1169 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_117 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_116_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_1177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_1179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_1186 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_116_1193 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_1203 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_116_1207 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_121 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_116_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_116_125 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_116_1261 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_116_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_1281 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_116_1284 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_129 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_116_1300 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_116_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_116_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_1331 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_1333 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_1336 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_116_1367 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_116_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_116_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_116_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_116_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_1461 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_1464 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_116_1472 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_116_1504 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_116_1520 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_1524 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_116_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_116_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_116_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_116_158 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_182 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_189 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_191 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_194 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_116_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_202 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_116_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_214 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_218 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_226 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_234 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_116_238 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_116_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_116_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_116_258 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_262 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_266 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_274 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_116_278 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_116_294 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_302 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_304 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_307 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_116_315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_116_324 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_328 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_330 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_333 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_341 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_116_345 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_116_353 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_359 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_366 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_116_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_116_370 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_116_386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_116_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_116_424 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_432 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_440 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_453 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_116_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_469 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_116_478 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_484 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_116_515 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_116_525 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_529 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_116_53 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_116_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_116_550 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_558 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_565 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_116_569 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_573 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_580 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_590 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_594 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_616 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_116_620 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_636 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_639 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_643 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_655 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_116_665 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_116_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_116_708 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_116_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_721 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_116_725 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_116_741 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_116_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_116_779 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_785 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_788 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_792 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_796 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_808 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_116_812 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_116_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_850 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_116_853 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_116_861 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_867 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_871 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_116_88 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_116_883 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_893 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_116_901 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_907 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_911 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_116_928 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_116_944 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_116_952 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_956 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_116_96 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_964 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_975 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_116_979 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_116_995 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_1014 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_1027 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_1035 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_117_1043 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_1059 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_1063 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_117_1070 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_1134 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_117_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_1142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_1146 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_117_1150 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_118 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_117_1182 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_1188 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_1200 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_1204 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_117_1212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_117_122 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_117_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_117_1252 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_1258 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_1266 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_117_1274 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_128 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_117_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_1284 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_117_1287 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_1297 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_1301 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_117_1311 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_1319 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_117_1322 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_117_1338 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_1346 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_117_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_1392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_1400 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_117_1404 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_1424 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_1427 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_117_1436 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_1468 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_1471 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_117_1479 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_117_1487 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_117_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_153 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_117_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_117_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_157 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_159 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_162 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_164 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_167 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_178 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_117_195 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_117_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_205 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_117_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_117_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_223 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_225 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_117_228 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_260 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_264 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_289 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_117_293 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_117_309 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_313 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_117_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_117_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_117_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_353 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_117_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_117_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_117_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_432 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_434 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_441 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_475 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_479 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_117_483 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_491 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_493 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_117_50 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_117_511 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_517 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_117_525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_117_541 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_553 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_557 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_117_561 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_565 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_117_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_117_58 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_117_586 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_590 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_117_594 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_117_606 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_117_622 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_630 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_117_64 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_652 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_654 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_117_657 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_117_665 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_671 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_117_674 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_68 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_117_706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_117_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_117_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_117_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_760 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_117_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_117_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_117_791 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_795 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_798 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_802 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_117_810 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_844 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_117_861 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_869 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_117_873 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_117_89 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_117_905 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_117_913 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_917 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_920 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_117_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_93 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_95 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_117_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_117_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_100 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_1001 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_1016 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_118_1020 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_118_1034 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_1042 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_118_1045 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_118_1077 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_118_1093 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_1097 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_118_1106 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_118_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_118_1130 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_1134 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_1137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_1141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_118_1151 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_1160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_1162 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_118_1165 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_1169 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_1175 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_118_1205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_122 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_1256 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_118_126 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_1264 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_118_1268 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_1276 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_1279 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_118_1283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_130 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_1301 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_118_1305 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_1317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_1320 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_118_1335 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_118_1367 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_1375 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_1398 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_1402 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_1406 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_118_1410 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_118_1444 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_1452 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_118_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_118_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_118_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_118_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_118_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_164 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_168 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_118_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_118_203 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_207 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_214 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_118_218 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_118_226 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_230 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_234 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_118_238 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_246 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_118_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_118_266 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_275 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_118_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_118_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_118_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_118_337 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_341 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_343 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_118_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_118_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_118_382 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_118_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_396 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_398 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_405 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_118_409 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_118_427 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_443 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_466 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_118_470 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_474 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_477 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_481 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_118_520 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_528 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_118_541 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_118_573 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_581 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_584 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_600 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_615 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_118_625 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_633 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_636 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_640 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_118_655 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_118_663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_688 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_118_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_118_692 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_118_708 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_118_716 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_720 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_722 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_118_725 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_729 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_118_733 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_118_741 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_118_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_751 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_118_759 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_118_767 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_771 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_775 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_782 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_118_786 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_118_802 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_118_810 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_814 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_118_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_834 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_836 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_118_846 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_85 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_850 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_852 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_118_855 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_87 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_118_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_118_921 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_118_928 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_932 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_118_936 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_952 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_954 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_96 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_966 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_970 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_118_974 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_118_982 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_986 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_990 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_994 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_119_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_119_1036 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_1040 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_1048 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_1070 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_1074 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_119_1084 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_119_1092 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_1104 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_1116 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_1120 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_1124 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_119_1128 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_1132 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_1150 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_1163 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_1167 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_1171 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_119_1175 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_1195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_1199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_119_1203 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_119_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_119_1217 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_1227 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_1229 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_1232 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_1251 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_1255 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_119_1259 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_1275 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_119_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_119_1316 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_119_1332 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_119_1340 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_1353 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_1360 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_119_1364 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_119_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_119_1372 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_1376 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_1399 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_1403 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_119_1407 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_119_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_119_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_1432 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_119_1439 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_1443 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_119_1452 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_119_1484 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_1488 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_119_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_119_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_119_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_195 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_119_199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_119_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_203 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_207 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_211 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_219 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_225 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_232 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_240 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_119_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_248 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_257 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_119_261 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_119_277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_281 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_119_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_119_302 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_310 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_319 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_119_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_119_360 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_376 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_388 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_119_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_408 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_412 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_431 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_435 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_119_439 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_119_447 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_453 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_467 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_475 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_477 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_119_490 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_119_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_119_50 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_507 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_517 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_519 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_119_533 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_537 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_540 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_549 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_555 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_119_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_119_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_574 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_578 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_58 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_119_588 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_622 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_626 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_119_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_119_67 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_714 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_119_721 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_119_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_731 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_119_762 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_766 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_769 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_119_777 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_119_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_119_791 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_795 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_798 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_119_808 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_119_840 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_119_848 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_119_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_119_864 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_874 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_878 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_888 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_119_892 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_910 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_928 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_119_932 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_119_942 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_119_950 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_954 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_962 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_119_966 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_978 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_119_982 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_119_990 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_119_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_11_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_11_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_11_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_11_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_11_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_11_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_11_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_11_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_11_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_11_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_11_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_11_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_11_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_11_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_11_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_11_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_11_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_11_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_11_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_11_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_11_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_11_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_11_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_120_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_120_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_120_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_1043 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_1046 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_1050 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_1062 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_120_1066 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_120_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_120_1082 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_120_1090 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_1094 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_1096 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_1117 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_1121 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_120_1125 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_120_1133 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_120_1139 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_120_1155 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_1159 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_1224 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_1226 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_1239 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_120_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_120_1276 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_1282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_120_1285 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_120_1301 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_1309 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_1326 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_1330 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_120_1334 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_1350 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_120_1353 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_120_1369 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_120_1377 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_1381 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_120_1389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_1397 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_140 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_120_1404 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_120_1420 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_1424 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_1426 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_1429 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_1433 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_1442 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_120_145 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_1452 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_120_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_120_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_120_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_120_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_120_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_120_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_120_195 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_120_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_120_203 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_207 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_210 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_217 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_223 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_234 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_238 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_120_242 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_246 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_120_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_266 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_269 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_120_277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_120_309 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_120_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_120_337 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_345 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_120_348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_120_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_120_380 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_388 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_399 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_120_403 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_411 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_459 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_120_514 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_520 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_120_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_120_537 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_541 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_543 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_552 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_586 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_590 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_120_594 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_620 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_624 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_120_628 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_120_660 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_120_668 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_672 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_120_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_120_708 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_120_716 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_720 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_120_723 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_120_733 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_120_741 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_120_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_120_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_120_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_120_828 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_120_844 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_853 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_857 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_861 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_863 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_120_870 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_120_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_120_897 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_901 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_903 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_906 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_120_914 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_930 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_120_938 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_120_954 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_120_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_964 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_120_968 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_978 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_120_982 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_120_990 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_994 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_120_997 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_121_1003 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_121_1011 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_1015 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_1023 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_1027 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_121_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_121_1047 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_121_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_121_1055 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_1059 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_1061 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_121_1074 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_121_1106 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_121_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_1130 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_1132 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_1140 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_1147 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_1155 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_1161 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_1165 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_1169 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_121_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_1181 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_121_1185 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_121_1201 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_1205 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_121_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_121_121 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_1213 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_1217 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_1225 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_1245 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_121_1249 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_125 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_1257 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_1259 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_1262 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_121_1266 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_1276 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_1287 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_129 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_1291 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_1298 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_121_1302 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_1310 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_1342 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_1346 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_121_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_1366 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_121_1370 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_121_1378 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_1382 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_1384 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_121_1387 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_121_1395 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_1399 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_1402 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_121_1416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_121_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_1438 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_1441 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_1448 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_121_1452 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_121_1484 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_1488 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_121_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_153 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_121_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_121_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_121_157 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_121_173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_185 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_121_189 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_193 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_121_196 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_121_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_121_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_121_249 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_257 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_121_260 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_121_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_121_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_121_364 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_121_380 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_121_388 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_394 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_401 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_121_405 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_121_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_442 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_446 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_121_450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_458 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_121_461 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_477 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_482 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_121_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_508 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_121_512 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_121_528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_121_536 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_540 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_542 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_555 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_121_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_576 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_121_580 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_584 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_588 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_121_592 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_121_624 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_121_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_636 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_121_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_649 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_652 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_656 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_121_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_121_668 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_672 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_674 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_677 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_684 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_121_688 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_121_704 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_708 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_121_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_121_728 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_121_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_121_736 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_742 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_121_745 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_761 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_121_764 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_121_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_121_791 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_795 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_797 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_800 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_810 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_814 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_826 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_834 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_838 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_846 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_848 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_121_862 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_876 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_121_880 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_121_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_920 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_121_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_929 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_937 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_941 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_121_945 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_961 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_121_965 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_969 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_121_972 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_988 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_990 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_100 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_1000 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_1003 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_1007 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_122_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_122_1025 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_122_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_1046 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_122_1050 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_122_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_1088 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_122_1092 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_122_1105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_122_1113 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_1117 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_122_1121 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_122_1137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_1156 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_1160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_1164 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_1168 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_122_1176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_1180 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_122_1183 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_1197 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_122_1201 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_122_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_1213 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_1215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_1218 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_1228 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_122_1232 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_1240 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_1248 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_1262 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_1274 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_1282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_1284 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_122_129 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_122_1291 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_1295 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_1304 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_1322 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_1326 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_1328 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_1331 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_122_1343 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_122_1355 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_122_1371 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_122_1402 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_1406 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_1409 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_122_1417 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_122_1449 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_1453 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_122_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_122_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_122_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_122_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_122_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_162 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_122_166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_186 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_188 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_194 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_122_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_228 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_232 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_236 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_238 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_122_258 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_264 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_272 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_292 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_122_296 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_122_312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_316 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_324 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_122_332 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_342 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_362 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_122_366 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_122_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_122_374 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_122_380 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_388 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_399 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_122_403 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_431 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_122_435 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_439 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_442 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_450 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_122_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_458 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_122_470 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_122_503 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_507 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_520 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_122_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_528 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_536 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_574 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_586 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_594 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_122_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_122_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_637 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_639 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_642 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_646 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_122_658 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_122_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_680 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_684 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_122_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_694 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_122_698 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_122_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_122_725 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_122_733 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_762 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_122_77 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_122_773 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_777 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_122_787 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_122_803 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_81 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_122_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_83 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_848 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_122_852 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_860 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_864 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_122_868 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_884 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_122_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_905 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_96 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_963 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_122_994 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_998 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_1000 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_1003 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_123_1011 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_123_1043 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_123_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_1059 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_1061 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_1078 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_123_1082 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_1086 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_1098 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_123_1106 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_1110 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_1119 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_1127 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_123_1141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_1145 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_1152 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_1183 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_1187 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_1189 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_1196 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_123_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_123_121 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_1215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_1229 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_1243 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_123_1247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_123_1255 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_1259 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_1261 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_123_1264 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_1272 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_1276 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_123_131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_1331 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_123_1339 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_1347 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_1359 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_1363 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_123_1367 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_123_1399 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_1407 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_1429 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_123_1433 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_1437 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_1439 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_123_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_123_1446 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_123_1478 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_123_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_123_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_123_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_123_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_123_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_184 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_123_188 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_192 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_123_196 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_123_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_123_204 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_123_224 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_257 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_123_261 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_123_277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_293 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_123_297 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_123_313 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_329 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_337 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_123_341 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_123_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_353 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_359 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_362 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_366 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_378 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_123_386 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_418 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_458 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_123_462 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_123_470 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_474 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_481 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_123_485 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_508 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_123_541 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_545 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_548 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_552 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_123_560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_123_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_574 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_578 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_123_582 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_586 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_590 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_123_594 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_604 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_607 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_611 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_621 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_123_625 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_123_633 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_637 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_123_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_123_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_123_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_123_689 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_123_697 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_701 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_123_721 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_123_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_123_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_123_745 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_751 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_760 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_764 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_123_768 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_123_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_123_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_793 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_800 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_123_804 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_820 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_824 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_832 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_123_840 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_123_848 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_123_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_123_862 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_868 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_123_876 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_123_892 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_123_900 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_904 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_123_908 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_916 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_123_919 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_932 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_123_940 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_972 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_980 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_123_984 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_992 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_123_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_124_1004 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_1008 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_124_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_1016 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_124_1020 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_124_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_1040 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_124_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_124_1076 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_124_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_1084 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_124_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_1097 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_124_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_1106 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_1120 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_1149 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_1163 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_124_1167 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_1187 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_1199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_124_1203 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_124_1219 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_1227 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_1231 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_124_1235 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_1239 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_124_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_1260 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_1272 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_1276 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_1278 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_124_1281 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_1290 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_1294 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_1298 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_124_1302 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_1310 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_124_1319 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_124_1335 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_124_1343 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_1347 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_1358 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_1360 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_124_1373 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_1381 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_124_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_124_1418 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_124_1434 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_1438 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_1440 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_1443 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_124_1451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_124_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_124_146 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_124_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_124_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_124_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_124_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_124_162 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_124_170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_124_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_183 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_185 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_124_188 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_124_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_124_220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_226 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_236 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_124_240 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_124_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_284 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_287 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_294 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_124_298 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_124_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_124_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_124_331 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_124_363 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_124_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_124_371 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_375 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_377 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_124_380 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_388 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_124_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_124_408 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_412 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_124_434 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_440 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_124_444 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_452 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_465 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_472 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_479 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_124_483 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_491 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_509 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_124_516 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_526 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_530 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_541 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_545 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_124_549 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_124_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_124_594 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_124_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_124_621 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_627 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_124_639 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_671 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_124_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_692 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_696 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_124_704 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_124_736 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_124_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_124_755 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_759 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_124_762 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_124_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_124_804 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_124_812 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_124_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_124_826 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_830 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_124_834 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_871 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_875 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_124_879 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_124_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_897 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_899 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_124_906 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_910 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_917 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_124_927 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_931 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_124_934 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_124_950 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_124_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_964 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_124_974 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_984 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_124_988 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_125_1012 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_1020 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_1023 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_1027 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_1037 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_125_1045 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_125_1061 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_125_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_125_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_125_1075 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_1089 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_125_1107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_1111 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_1121 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_1129 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_1133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_1144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_1148 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_125_115 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_125_1152 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_1160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_1163 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_125_1167 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_1171 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_1180 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_1187 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_119 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_1191 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_125_1195 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_125_1203 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_125_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_1213 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_1217 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_125_122 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_125_1225 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_125_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_1249 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_1252 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_125_1260 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_1276 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_128 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_1289 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_1297 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_125_1301 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_1309 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_1311 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_1317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_1331 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_125_1335 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_125_1343 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_1347 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_125_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_1355 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_1357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_125_1360 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_1368 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_1370 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_125_1377 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_125_138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_125_1393 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_1403 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_125_1407 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_125_1413 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_1417 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_125_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_125_1438 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_1444 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_1448 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_125_1462 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_125_1478 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_125_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_125_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_125_151 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_125_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_125_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_125_167 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_186 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_194 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_125_198 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_125_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_125_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_210 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_125_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_225 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_233 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_125_237 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_125_253 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_257 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_264 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_268 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_125_272 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_125_280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_125_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_125_302 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_310 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_125_364 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_125_396 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_125_412 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_125_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_435 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_439 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_125_443 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_125_459 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_125_467 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_471 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_125_474 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_125_490 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_494 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_125_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_507 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_125_511 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_125_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_125_535 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_539 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_125_543 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_551 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_125_560 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_125_577 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_125_609 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_125_625 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_125_633 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_637 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_125_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_125_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_715 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_125_725 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_125_757 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_763 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_770 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_125_786 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_125_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_125_826 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_832 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_125_840 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_125_848 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_856 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_125_859 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_863 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_866 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_87 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_125_874 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_125_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_888 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_125_896 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_900 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_125_908 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_125_91 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_938 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_125_942 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_125_950 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_954 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_961 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_125_969 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_973 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_976 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_125_980 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_125_988 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_992 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_125_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_1001 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_126_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_1016 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_1020 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_1034 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_1036 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_126_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_126_1047 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_1051 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_1058 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_1062 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_1066 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_126_1070 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_126_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_1086 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_126_1089 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_1097 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_126_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_1118 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_112 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_1120 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_126_1123 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_1142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_126_1146 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_126_1156 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_1176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_126_1180 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_1184 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_1186 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_126_1189 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_1193 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_1195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_1198 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_120 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_1210 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_1218 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_1228 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_1232 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_126_1236 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_126_124 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_1240 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_1274 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_1289 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_1293 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_126_1297 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_1301 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_1330 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_1338 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_126_1342 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_1346 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_1354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_126_1362 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_1368 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_126_1372 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_126_1380 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_126_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_1390 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_1392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_1399 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_1403 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_1413 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_1420 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_126_1424 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_126_1440 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_126_1448 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_1452 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_126_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_126_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_126_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_126_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_126_157 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_126_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_126_173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_126_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_183 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_185 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_188 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_190 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_193 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_126_197 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_126_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_126_205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_211 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_126_214 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_246 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_126_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_254 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_262 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_270 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_278 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_292 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_126_296 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_126_312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_316 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_126_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_325 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_327 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_126_330 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_126_338 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_126_348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_126_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_380 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_126_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_388 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_126_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_408 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_429 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_126_442 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_448 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_126_452 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_126_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_469 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_479 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_483 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_126_487 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_126_503 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_126_511 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_515 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_537 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_126_541 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_126_557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_565 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_126_569 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_126_577 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_581 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_584 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_126_592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_600 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_126_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_126_637 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_126_653 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_661 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_665 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_684 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_126_688 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_126_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_126_720 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_730 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_126_734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_126_754 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_126_77 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_126_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_804 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_81 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_126_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_126_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_822 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_824 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_830 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_834 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_836 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_126_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_857 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_126_865 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_126_881 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_885 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_89 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_126_892 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_126_926 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_126_93 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_126_963 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_997 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_1006 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_1010 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_1012 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_1021 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_127_103 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_1035 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_1043 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_1046 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_1054 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_1058 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_1083 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_127_1091 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_127_1123 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_127_1147 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_127_1159 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_127_1175 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_1183 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_1187 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_1191 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_127_1195 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_1203 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_1212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_1219 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_1229 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_127_1233 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_1265 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_1283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_1287 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_1293 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_1297 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_1299 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_127_1302 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_1318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_1320 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_1327 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_1335 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_127_1339 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_1347 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_1355 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_1357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_1366 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_1374 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_127_1378 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_1390 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_1393 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_1399 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_127_1407 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_127_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_127_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_127_156 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_127_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_127_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_180 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_189 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_193 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_197 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_127_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_201 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_218 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_232 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_127_236 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_252 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_260 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_264 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_268 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_127_272 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_293 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_127_297 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_313 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_328 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_342 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_344 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_127_347 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_127_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_373 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_375 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_382 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_390 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_127_394 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_410 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_414 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_127_417 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_430 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_433 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_437 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_441 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_127_444 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_452 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_127_455 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_127_487 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_495 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_127_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_127_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_547 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_551 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_555 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_573 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_127_577 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_585 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_589 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_593 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_607 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_127_611 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_619 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_623 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_631 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_635 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_671 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_127_675 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_707 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_716 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_719 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_726 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_127_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_127_730 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_127_746 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_754 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_760 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_767 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_127_771 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_779 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_786 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_796 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_800 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_127_804 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_127_820 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_828 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_832 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_835 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_127_839 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_856 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_127_859 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_875 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_879 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_887 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_89 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_897 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_901 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_905 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_911 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_127_915 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_929 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_932 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_936 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_942 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_946 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_958 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_966 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_97 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_970 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_127_974 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_990 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_1006 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_1010 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_1014 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_1016 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_1025 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_128_1034 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_1050 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_1054 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_1057 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_1068 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_1072 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_1076 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_128_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_128_1091 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_1111 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_1115 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_1119 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_1123 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_1145 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_1149 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_1153 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_1176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_1189 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_1197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_1201 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_1205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_1211 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_1214 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_1218 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_1220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_128_1227 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_1235 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_1239 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_124 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_128_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_128_1260 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_1268 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_128_1274 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_1306 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_1322 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_1330 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_1337 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_1345 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_1349 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_128_1353 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_1363 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_1377 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_1381 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_1389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_1420 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_128_1424 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_128_1440 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_1448 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_1452 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_128_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_128_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_128_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_182 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_188 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_196 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_198 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_128_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_201 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_216 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_230 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_234 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_238 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_242 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_246 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_252 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_259 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_128_269 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_128_301 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_327 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_335 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_345 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_128_356 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_128_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_128_372 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_128_402 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_434 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_436 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_439 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_443 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_453 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_128_472 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_128_504 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_128_514 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_530 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_128_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_566 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_573 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_128_584 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_600 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_128_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_128_621 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_629 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_635 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_639 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_646 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_648 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_657 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_661 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_665 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_128_685 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_128_701 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_713 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_723 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_727 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_128_731 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_739 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_743 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_128_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_128_825 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_857 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_861 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_865 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_873 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_881 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_883 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_898 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_902 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_904 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_907 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_911 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_928 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_932 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_128_944 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_952 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_956 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_128_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_128_976 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_984 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_988 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_994 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_128_998 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_1000 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_1003 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_129_1007 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_129_1015 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_129_1021 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_129_1037 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_129_1045 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_1049 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_129_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_1051 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_1054 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_1058 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_1062 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_129_1070 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_129_1086 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_129_1094 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_1098 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_1108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_129_1115 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_1125 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_1133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_1140 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_1153 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_1160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_1164 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_1168 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_1172 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_129_1184 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_1188 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_1191 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_129_1195 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_129_1203 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_129_121 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_1212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_1216 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_1220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_1233 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_129_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_129_1253 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_129_1261 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_1265 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_1267 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_1270 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_129_1274 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_129 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_1290 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_1294 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_129_1298 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_129_1314 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_129_1324 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_1328 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_129_1332 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_1364 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_1371 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_1375 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_129_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_129_1399 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_129_1413 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_1417 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_129_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_129_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_129_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_129_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_129_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_129_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_129_160 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_129_168 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_178 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_129_182 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_198 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_129_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_200 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_129_203 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_207 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_218 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_227 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_238 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_248 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_129_252 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_129_268 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_272 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_275 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_293 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_129_297 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_129_313 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_319 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_129_322 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_129_330 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_129_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_129_373 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_129_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_129_388 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_129_396 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_129_412 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_420 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_435 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_437 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_129_440 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_129_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_464 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_470 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_129_474 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_129_490 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_494 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_512 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_522 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_526 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_129_530 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_129_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_566 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_129_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_129_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_129_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_129_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_129_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_129_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_129_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_129_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_129_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_129_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_861 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_865 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_869 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_893 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_900 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_914 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_129_932 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_129_940 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_944 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_946 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_949 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_129_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_961 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_964 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_977 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_981 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_129_985 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_129_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_12_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_12_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_12_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_12_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_12_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_12_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_12_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_12_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_12_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_12_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_12_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_12_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_12_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_12_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_12_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_12_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_12_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_12_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_12_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_12_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_12_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_12_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_12_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_12_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_1005 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_130_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_1019 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_1026 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_1034 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_130_1038 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_1048 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_1056 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_1078 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_130_1082 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_1098 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_130_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_1106 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_1110 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_1114 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_130_1118 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_130_1134 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_1141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_130_115 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_130_1151 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_130_1167 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_130_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_1181 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_1183 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_130_1186 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_119 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_130_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_1208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_1212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_1216 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_1229 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_130_1233 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_1250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_130_1254 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_1258 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_1268 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_130_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_1294 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_1298 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_130_1302 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_1322 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_130_1326 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_130_1336 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_130_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_130_1358 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_1362 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_1376 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_130_1389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_1453 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_130_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_130_150 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_130_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_130_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_130_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_130_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_130_158 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_162 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_165 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_185 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_189 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_130_193 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_130_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_130_210 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_130_220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_224 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_226 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_130_229 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_240 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_130_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_130_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_130_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_130_298 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_306 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_310 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_327 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_130_331 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_130_343 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_130_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_130_375 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_130_383 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_130_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_130_424 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_130_438 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_448 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_130_452 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_130_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_130_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_130_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_538 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_540 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_543 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_130_553 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_130_585 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_601 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_130_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_609 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_611 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_614 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_625 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_130_629 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_130_645 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_649 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_652 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_656 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_660 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_130_679 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_130_695 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_703 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_130_708 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_130_724 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_130_732 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_736 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_130_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_130_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_785 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_130_789 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_793 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_797 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_130_805 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_813 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_820 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_823 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_831 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_833 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_836 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_130_844 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_130_860 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_868 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_130_871 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_879 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_881 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_884 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_892 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_896 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_900 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_904 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_908 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_130_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_130_944 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_130_952 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_956 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_130_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_968 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_970 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_130_973 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_130_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_995 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_998 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_1000 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_1002 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_1005 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_131_1009 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_131_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_131_1023 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_131_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_1043 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_1046 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_1050 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_131_1061 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_1070 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_131_1074 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_131_1090 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_131_1098 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_131_1106 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_1110 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_1112 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_1125 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_131_1129 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_113 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_1133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_131_1151 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_131_1167 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_117 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_1177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_1184 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_1196 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_131_1200 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_1204 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_121 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_1211 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_1214 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_1225 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_131_1229 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_1239 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_1242 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_1249 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_131_1253 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_131_1261 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_1265 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_1267 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_131_1270 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_128 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_1283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_1287 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_131_1291 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_131_1307 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_1311 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_1325 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_131_1332 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_131_1342 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_131_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_1365 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_131_1380 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_140 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_131_1412 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_131_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_131_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_148 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_131_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_131_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_151 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_155 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_131_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_131_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_162 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_180 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_131_184 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_188 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_190 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_193 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_131_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_202 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_131_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_218 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_230 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_234 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_131_238 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_131_254 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_262 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_131_269 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_131_277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_281 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_131_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_131_302 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_316 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_131_324 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_334 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_131_338 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_131_372 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_131_388 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_399 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_131_403 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_407 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_409 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_131_420 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_424 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_131_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_131_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_131_476 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_480 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_131_484 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_131_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_131_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_131_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_539 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_541 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_131_544 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_131_560 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_581 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_585 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_131_589 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_593 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_131_596 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_131_628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_636 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_131_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_131_657 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_131_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_677 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_131_681 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_689 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_692 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_704 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_706 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_719 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_723 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_131_727 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_131_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_731 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_733 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_736 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_758 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_131_762 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_778 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_131_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_791 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_795 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_808 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_812 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_816 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_820 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_131_824 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_131_840 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_848 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_867 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_871 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_875 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_879 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_131_883 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_899 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_902 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_131_906 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_921 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_131_928 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_131_944 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_131_952 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_956 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_958 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_961 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_971 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_981 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_131_985 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_131_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_132_1003 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_132_1009 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_132_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_132_1019 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_1027 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_132_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_1046 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_132_1050 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_1058 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_132_1063 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_132_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_1106 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_132_1114 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_132_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_1126 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_1132 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_1146 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_1148 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_1155 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_132_1159 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_1167 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_132_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_132_1183 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_132_1215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_1225 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_132_1235 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_1239 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_132_124 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_132_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_132_1260 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_1268 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_1275 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_1279 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_132_1283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_132_1299 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_132_130 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_132_1307 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_1311 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_132_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_1319 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_1325 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_1339 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_1345 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_132_1349 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_1355 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_1361 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_132_1371 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_132_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_132_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_132_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_132_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_132_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_132_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_132_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_132_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_162 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_164 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_132_170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_193 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_132_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_132_207 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_213 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_132_222 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_228 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_238 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_242 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_132_261 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_267 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_271 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_132_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_290 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_297 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_132_301 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_305 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_309 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_313 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_326 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_330 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_132_334 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_342 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_132_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_132_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_132_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_388 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_132_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_132_424 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_132_432 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_436 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_132_439 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_132_455 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_459 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_132_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_132_482 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_488 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_132_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_132_500 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_132_516 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_132_525 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_536 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_542 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_549 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_132_553 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_132_569 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_132_577 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_581 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_585 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_594 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_132_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_609 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_615 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_132_619 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_651 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_654 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_132_662 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_670 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_132_683 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_132_699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_132_706 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_714 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_718 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_725 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_132_733 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_760 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_132_764 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_132_798 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_814 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_132_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_858 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_862 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_132_866 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_132_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_895 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_899 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_906 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_910 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_914 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_132_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_132_931 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_132_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_955 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_132_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_966 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_979 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_983 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_132_987 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_1007 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_133_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_133_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_1048 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_1054 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_133_1058 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_1062 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_133_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_1075 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_1077 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_133_1080 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_1089 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_1104 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_1116 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_133_1123 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_133_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_1145 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_133_1149 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_133_1165 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_1175 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_133_1178 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_1186 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_1196 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_133_1200 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_1204 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_133_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_1219 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_1235 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_133_1239 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_1255 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_1257 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_1260 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_1264 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_1276 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_1289 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_133_1293 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_133_1309 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_1319 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_1331 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_1341 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_133_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_1359 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_133_1363 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_133_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_133_1395 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_133_1411 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_133_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_133_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_133_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_133_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_133_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_133_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_133_178 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_186 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_190 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_194 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_133_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_201 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_218 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_223 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_227 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_133_257 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_263 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_133_267 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_133_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_290 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_292 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_305 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_319 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_323 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_325 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_133_328 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_336 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_133_347 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_133_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_133_365 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_369 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_371 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_380 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_390 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_133_394 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_133_410 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_133_418 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_133_437 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_441 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_448 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_133_452 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_505 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_133_509 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_133_541 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_133_549 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_553 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_565 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_133_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_133_586 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_133_596 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_606 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_610 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_620 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_133_624 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_133_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_133_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_645 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_647 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_650 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_133_658 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_133_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_690 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_694 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_698 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_715 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_133_719 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_723 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_133_727 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_133_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_735 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_748 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_760 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_133_764 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_133_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_133_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_133_796 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_802 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_133_806 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_133_822 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_832 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_133_836 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_840 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_849 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_133_857 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_873 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_875 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_894 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_902 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_910 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_928 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_133_932 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_936 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_938 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_941 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_133_949 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_961 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_971 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_981 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_985 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_133_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_999 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_1002 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_1004 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_134_1007 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_134_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_1015 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_134_1019 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_1027 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_134_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_1041 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_134_1045 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_1055 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_1065 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_1071 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_134_1075 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_1079 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_134_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_1088 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_1092 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_1105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_1107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_134_1118 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_134_1150 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_1176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_1188 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_1200 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_1204 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_134_1208 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_134_1214 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_1218 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_1220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_1231 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_1235 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_1239 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_134_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_1252 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_1254 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_134_1257 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_134_1265 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_1269 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_134_1290 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_134_1306 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_1323 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_1337 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_134_1341 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_134_1373 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_1381 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_134_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_134_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_134_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_134_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_134_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_134_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_134_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_134_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_134_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_134_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_134_211 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_134_219 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_225 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_229 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_239 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_261 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_271 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_134_275 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_307 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_134_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_325 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_327 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_330 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_338 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_134_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_134_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_134_378 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_134_386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_134_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_424 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_427 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_134_441 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_447 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_134_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_459 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_134_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_134_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_134_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_134_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_134_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_611 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_134_619 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_134_627 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_631 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_642 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_655 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_134_659 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_134_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_671 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_134_679 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_134_695 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_701 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_704 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_708 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_718 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_134_722 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_134_738 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_134_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_756 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_134_760 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_134_792 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_800 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_802 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_809 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_813 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_820 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_823 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_830 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_134_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_856 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_860 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_864 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_134_868 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_884 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_134_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_893 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_896 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_900 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_904 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_908 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_134_916 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_134_948 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_956 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_963 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_967 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_969 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_978 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_982 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_986 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_134_990 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_134_998 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_1005 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_1012 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_1016 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_135_1020 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_1030 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_1033 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_1041 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_1053 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_135_1057 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_135_106 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_135_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_135_1083 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_1089 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_1092 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_1096 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_1107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_1111 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_1115 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_1127 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_135_1147 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_1161 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_1171 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_135_1175 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_1179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_1190 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_1194 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_135_1198 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_1212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_1222 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_1224 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_1235 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_1247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_1251 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_1255 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_1265 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_135_1269 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_1283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_135_1287 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_135_1319 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_135_1335 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_135_1343 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_1347 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_135_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_135_138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_135_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_135_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_135_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_135_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_135_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_135_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_135_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_135_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_135_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_135_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_231 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_235 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_239 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_135_248 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_135_256 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_260 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_135_263 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_135_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_135_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_135_302 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_306 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_320 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_135_324 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_135_340 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_135_348 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_135_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_135_373 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_377 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_382 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_135_396 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_135_412 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_420 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_430 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_442 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_446 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_450 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_135_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_135_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_494 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_135_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_135_507 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_511 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_513 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_516 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_526 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_135_530 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_135_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_566 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_135_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_135_586 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_135_594 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_601 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_135_609 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_135_625 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_135_633 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_637 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_135_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_649 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_652 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_656 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_135_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_660 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_675 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_678 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_690 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_135_694 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_724 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_135_728 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_135_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_135_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_748 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_135_751 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_767 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_135_771 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_779 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_135_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_135_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_819 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_821 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_824 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_834 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_135_838 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_135_844 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_135_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_135_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_135_89 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_894 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_897 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_135_905 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_135_913 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_917 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_920 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_135_928 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_93 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_135_936 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_940 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_944 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_948 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_95 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_970 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_135_974 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_135_980 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_988 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_990 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_136_1008 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_136_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_136_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_1035 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_1045 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_1057 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_1061 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_136_1065 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_136_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_1097 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_136_1105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_136_1137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_1153 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_136_1167 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_1176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_1180 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_136_1184 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_1188 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_136_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_136_1208 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_136_1216 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_1220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_1227 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_136_1231 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_136_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_136_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_1260 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_1267 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_136_1271 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_136_1303 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_1311 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_136_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_136_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_136_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_136_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_136_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_136_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_136_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_136_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_136_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_136_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_136_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_136_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_136_211 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_235 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_136_239 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_136_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_136_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_136_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_136_353 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_369 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_136_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_371 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_388 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_136_395 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_136_429 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_136_437 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_441 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_136_444 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_136_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_544 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_548 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_136_552 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_136_568 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_580 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_584 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_586 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_136_589 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_136_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_601 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_136_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_637 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_136_640 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_136_648 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_652 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_136_656 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_672 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_136_679 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_743 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_136_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_136_755 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_767 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_774 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_778 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_136_782 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_790 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_793 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_803 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_136_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_136_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_136_834 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_136_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_846 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_849 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_859 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_863 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_136_867 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_136_883 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_136_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_136_897 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_901 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_904 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_908 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_920 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_932 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_936 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_136_940 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_136_948 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_952 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_954 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_967 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_136_975 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_136_991 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_999 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_1007 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_137_1011 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_137_1027 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_1037 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_1041 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_1045 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_1057 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_137_1061 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_137_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_137_1083 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_1091 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_1094 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_1104 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_1111 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_137_1115 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_1119 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_137_1123 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_137_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_137_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_137_1146 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_1150 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_1161 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_137_1165 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_137_1171 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_137_1203 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_137_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_1213 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_1216 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_1226 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_1230 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_137_1234 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_137_1266 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_137_1274 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_1310 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_1314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_1318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_137_1322 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_137_1338 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_1346 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_137_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_137_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_137_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_137_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_137_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_137_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_137_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_137_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_137_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_137_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_137_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_137_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_137_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_137_255 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_137_271 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_137_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_137_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_137_302 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_310 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_137_325 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_333 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_337 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_137_347 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_351 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_137_370 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_374 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_382 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_137_386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_137_402 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_410 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_137_413 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_137_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_444 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_447 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_449 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_452 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_137_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_137_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_506 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_510 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_137_514 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_137_546 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_137_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_566 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_137_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_576 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_137_587 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_593 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_137_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_137_613 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_621 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_623 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_626 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_644 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_137_648 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_137_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_137_664 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_672 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_675 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_687 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_137_691 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_707 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_137_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_137_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_137_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_137_760 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_764 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_766 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_137_769 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_137_777 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_137_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_787 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_789 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_792 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_137_800 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_804 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_137_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_137_843 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_864 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_874 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_878 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_137_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_137_890 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_894 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_897 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_901 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_137_916 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_137_928 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_137_944 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_137_952 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_956 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_964 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_966 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_137_969 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_137_985 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_998 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_1002 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_1005 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_1009 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_138_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_1021 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_138_1025 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_138_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_138_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_1045 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_1062 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_1066 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_1070 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_1074 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_1078 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_138_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_1082 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_1111 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_1121 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_1129 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_138_1133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_1137 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_138_1143 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_1149 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_1163 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_138_1176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_1180 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_1182 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_1195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_1201 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_138_1205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_1213 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_1226 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_138_1247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_138_1263 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_1271 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_1274 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_1305 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_1311 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_1322 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_138_1326 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_138_1358 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_138_1374 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_1382 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_138_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_138_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_138_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_138_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_138_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_138_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_138_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_138_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_138_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_138_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_138_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_138_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_138_266 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_138_274 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_278 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_291 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_298 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_138_302 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_308 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_138_312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_316 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_138_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_138_353 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_361 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_364 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_138_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_374 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_138_378 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_138_386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_138_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_400 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_403 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_411 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_138_423 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_429 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_433 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_435 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_438 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_138_445 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_449 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_452 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_138_472 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_138_488 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_495 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_497 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_138_500 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_536 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_138_539 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_555 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_138_558 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_138_590 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_138_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_138_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_138_621 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_629 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_631 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_637 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_138_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_138_657 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_663 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_138_670 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_138_679 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_138_695 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_706 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_710 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_714 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_728 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_138_732 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_758 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_762 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_138_766 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_138_798 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_814 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_138_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_138_850 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_138_858 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_862 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_866 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_138_870 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_874 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_878 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_138_896 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_902 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_138_906 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_910 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_913 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_138_921 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_937 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_940 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_138_950 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_954 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_969 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_138_973 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_138_979 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_995 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_138_998 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_1005 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_139_1009 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_1013 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_1015 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_139_1018 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_1032 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_139_1036 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_1047 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_1051 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_139_1061 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_1074 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_139_1078 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_1084 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_1098 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_139_1113 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_139_1129 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_139_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_1154 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_1168 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_1172 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_139_1176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_1180 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_1184 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_139_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_139_1212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_1216 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_1219 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_1230 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_1240 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_1271 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_1275 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_139_1331 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_1347 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_139_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_139_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_139_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_139_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_139_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_139_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_139_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_139_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_139_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_139_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_139_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_139_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_139_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_139_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_139_294 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_316 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_320 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_328 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_139_332 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_338 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_342 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_139_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_139_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_139_365 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_369 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_371 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_139_374 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_139_390 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_139_398 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_402 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_404 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_407 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_409 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_412 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_420 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_424 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_139_435 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_441 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_139_493 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_537 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_139_541 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_545 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_139_554 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_139_560 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_581 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_585 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_139_589 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_593 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_601 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_139_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_637 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_139_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_657 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_659 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_139_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_662 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_139_677 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_139_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_139_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_789 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_139_793 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_139_801 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_805 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_813 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_139_817 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_139_833 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_837 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_840 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_850 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_139_857 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_139_873 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_139_881 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_885 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_888 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_900 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_907 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_911 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_139_915 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_919 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_139_928 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_932 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_936 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_139_940 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_946 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_950 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_964 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_968 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_972 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_976 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_978 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_981 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_985 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_13_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_13_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_13_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_13_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_13_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_13_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_13_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_13_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_13_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_13_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_13_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_13_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_13_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_13_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_13_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_13_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_13_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_13_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_13_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_13_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_13_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_13_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_13_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_1000 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_1007 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_140_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_1011 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_1015 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_1019 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_1023 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_1027 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_140_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_1037 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_1045 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_1049 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_1053 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_1063 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_1078 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_140_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_1086 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_1090 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_1094 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_1098 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_140_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_1114 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_140_1120 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_140_1136 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_140_1144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_1148 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_1155 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_1162 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_1180 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_1184 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_1186 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_140_1216 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_140_1222 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_1234 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_140_1238 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_140_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_1276 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_1279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_1287 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_140_1291 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_140_1305 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_140_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_140_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_140_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_140_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_140_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_140_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_140_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_140_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_140_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_140_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_140_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_140_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_140_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_140_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_140_266 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_274 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_306 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_323 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_334 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_342 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_140_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_366 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_140_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_140_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_394 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_397 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_405 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_140_417 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_427 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_439 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_447 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_140_455 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_459 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_470 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_472 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_479 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_140_483 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_140_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_503 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_140_510 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_514 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_525 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_529 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_140_537 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_553 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_556 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_558 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_140_588 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_140_596 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_600 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_140_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_140_621 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_629 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_140_633 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_140_665 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_140_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_140_708 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_720 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_140_724 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_140_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_140_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_140_763 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_140_771 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_775 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_778 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_785 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_140_789 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_140_805 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_813 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_824 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_828 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_140_832 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_140_848 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_140_856 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_860 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_862 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_876 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_880 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_884 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_140_896 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_900 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_913 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_140_917 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_921 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_924 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_140_934 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_946 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_948 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_967 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_971 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_975 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_979 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_981 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_988 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_992 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_140_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_1005 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_141_1019 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_1029 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_1033 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_1037 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_1054 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_1070 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_1072 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_1109 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_1113 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_141_1117 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_1121 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_1123 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_1130 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_1134 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_1145 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_1149 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_1153 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_1161 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_141_1171 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_1175 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_1183 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_1187 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_1191 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_1195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_1205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_1212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_1216 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_1224 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_1255 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_141_1259 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_1275 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_141_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_141_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_141_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_141_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_141_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_141_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_141_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_141_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_141_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_141_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_141_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_141_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_141_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_141_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_141_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_141_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_290 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_298 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_306 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_338 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_359 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_372 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_380 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_141_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_388 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_391 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_141_407 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_413 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_458 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_462 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_470 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_141_474 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_141_490 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_494 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_507 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_141_529 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_141_547 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_621 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_141_631 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_637 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_141_644 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_141_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_141_660 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_668 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_141_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_141_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_141_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_141_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_141_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_141_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_141_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_141_831 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_835 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_845 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_849 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_141_857 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_865 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_895 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_899 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_901 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_908 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_928 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_930 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_141_964 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_968 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_979 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_987 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_142_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_1019 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_1026 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_142_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_1041 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_1055 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_1061 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_1063 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_142_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_1093 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_1097 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_1105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_1111 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_1115 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_142_1119 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_1123 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_1132 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_1163 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_142_1167 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_1224 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_1228 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_142_1238 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_1247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_142_1251 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_142_1283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_142_1299 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_142_1307 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_1311 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_142_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_142_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_142_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_142_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_142_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_142_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_142_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_142_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_142_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_142_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_142_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_142_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_142_211 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_142_219 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_223 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_239 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_142_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_142_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_142_258 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_291 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_142_295 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_142_303 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_307 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_310 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_336 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_142_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_388 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_396 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_427 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_458 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_142_466 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_142_482 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_490 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_505 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_511 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_529 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_142_537 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_545 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_547 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_577 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_585 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_142_589 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_593 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_595 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_616 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_624 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_142_628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_662 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_671 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_142_679 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_142_695 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_706 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_727 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_731 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_735 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_758 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_142_762 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_142_794 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_142_810 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_814 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_142_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_142_850 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_142_858 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_862 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_876 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_884 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_893 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_902 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_910 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_142_941 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_945 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_142_954 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_975 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_983 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_987 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_1010 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_1016 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_143_1026 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_1037 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_1047 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_1057 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_1118 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_1126 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_1130 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_1134 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_143_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_143_1154 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_1158 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_1162 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_143_1174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_143_1190 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_1198 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_143_1212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_1222 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_1226 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_1228 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_143_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_143_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_143_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_143_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_143_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_143_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_143_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_143_1389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_143_1405 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_143_1413 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_1417 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_143_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_143_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_143_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_143_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_143_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_143_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_143_1572 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_143_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_143_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_143_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_231 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_143_289 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_297 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_343 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_143_351 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_372 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_376 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_407 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_423 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_143_431 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_449 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_461 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_143_469 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_473 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_480 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_488 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_506 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_533 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_551 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_143_573 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_143_589 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_143_627 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_143_635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_143_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_143_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_143_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_681 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_143_684 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_143_700 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_708 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_143_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_143_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_143_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_143_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_787 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_791 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_801 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_805 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_143_809 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_143_825 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_143_833 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_843 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_143_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_856 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_870 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_874 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_878 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_143_909 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_913 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_976 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_143_980 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_984 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_10 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_1009 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_1013 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_1026 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_103 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_1033 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_1049 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_1068 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_1084 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_111 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_1117 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_1119 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_1137 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_144_1141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_1153 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_1161 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_144_117 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_144_1177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_1185 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_1189 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_1197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_1203 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_1219 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_1227 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_1230 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_1232 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_1243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_1259 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_144_1262 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_1270 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_1274 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_144_1279 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_1287 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_1291 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_1294 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_1297 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_1316 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_1321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_1325 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_1329 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_1332 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_144_1347 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_1355 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_1363 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_1367 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_1371 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_1387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_1395 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_1399 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_14 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_1402 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_144_1407 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_144_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_1437 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_1441 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_144_1447 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_1455 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_144_1461 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_1469 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_144_147 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_144_1472 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_1480 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_1484 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_144_1489 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_1497 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_1503 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_144_1507 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_1523 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_144_1531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_1539 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_1542 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_144_1547 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_1563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_1567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_1573 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_1577 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_144_159 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_181 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_144_187 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_144_19 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_195 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_144_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_201 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_238 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_242 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_263 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_27 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_285 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_289 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_293 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_320 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_324 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_327 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_33 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_331 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_355 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_359 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_363 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_144_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_404 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_448 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_472 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_474 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_144_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_506 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_53 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_538 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_542 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_573 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_144_579 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_601 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_144_607 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_144_61 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_629 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_144_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_640 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_644 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_144_649 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_682 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_686 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_691 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_695 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_144_717 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_725 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_733 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_741 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_757 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_144_761 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_769 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_144_77 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_777 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_799 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_803 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_817 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_823 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_839 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_144_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_850 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_859 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_861 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_864 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_868 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_874 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_892 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_900 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_908 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_927 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_93 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_933 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_937 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_943 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_97 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_977 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_979 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_982 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_987 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_991 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_14_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_14_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_14_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_14_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_14_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_14_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_14_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_14_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_14_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_14_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_14_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_14_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_14_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_14_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_14_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_14_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_14_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_14_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_14_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_14_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_14_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_14_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_14_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_14_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_15_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_15_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_15_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_15_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_15_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_15_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_15_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_15_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_15_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_15_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_15_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_15_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_15_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_15_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_15_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_15_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_15_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_15_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_15_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_15_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_15_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_15_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_15_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_16_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_16_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_16_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_16_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_16_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_16_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_16_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_16_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_16_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_16_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_16_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_16_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_16_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_16_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_16_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_16_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_16_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_16_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_16_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_16_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_16_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_16_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_16_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_16_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_17_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_17_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_17_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_17_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_17_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_17_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_17_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_17_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_17_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_17_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_17_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_17_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_17_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_17_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_17_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_17_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_17_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_17_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_17_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_17_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_17_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_17_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_17_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_18_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_18_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_18_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_18_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_18_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_18_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_18_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_18_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_18_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_18_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_18_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_18_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_18_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_18_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_18_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_18_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_18_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_18_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_18_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_18_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_18_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_18_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_18_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_18_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_19_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_19_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_19_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_19_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_19_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_19_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_19_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_19_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_19_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_19_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_19_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_19_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_19_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_19_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_19_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_19_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_19_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_19_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_19_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_19_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_19_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_19_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_19_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_1005 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_1013 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_1047 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_1_1051 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_1059 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_1063 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_1074 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_1_1105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_1_1121 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_1129 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_1133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_1_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_1_1154 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_1162 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_1164 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_1194 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_1_1198 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_1_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_1217 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_1219 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_1222 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_1274 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_1287 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_1_1295 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_1_1327 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_1343 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_1347 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_1_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_1_1367 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_1375 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_1_1409 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_1417 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_1424 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_1431 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_1_1439 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_1_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_1_1471 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_1487 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_1_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_1_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_1_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_1_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_1_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_1_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_1_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_1_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_533 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_536 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_1_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_1_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_1_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_1_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_1_813 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_845 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_849 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_1_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_862 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_1_895 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_911 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_921 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_1_932 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_1_964 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_1_980 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_988 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_992 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_998 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_20_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_20_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_20_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_20_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_20_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_20_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_20_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_20_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_20_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_20_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_20_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_20_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_20_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_20_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_20_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_20_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_20_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_20_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_20_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_20_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_20_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_20_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_20_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_20_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_21_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_21_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_21_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_21_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_21_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_21_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_21_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_21_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_21_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_21_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_21_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_21_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_21_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_21_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_21_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_21_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_21_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_21_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_21_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_21_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_21_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_21_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_21_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_22_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_22_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_22_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_22_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_22_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_22_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_22_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_22_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_22_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_22_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_22_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_22_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_22_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_22_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_22_353 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_369 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_22_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_22_377 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_22_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_22_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_22_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_22_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_22_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_22_692 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_700 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_22_713 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_22_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_22_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_22_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_22_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_23_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_23_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_23_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_23_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_23_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_23_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_23_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_23_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_23_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_23_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_23_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_23_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_23_391 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_423 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_23_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_23_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_23_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_547 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_551 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_553 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_23_556 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_23_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_23_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_23_618 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_23_631 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_23_647 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_23_679 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_687 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_691 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_695 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_697 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_706 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_23_721 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_23_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_23_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_745 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_753 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_757 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_23_761 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_777 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_23_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_23_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_23_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_23_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_24_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_24_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_24_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_24_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_24_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_24_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_24_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_24_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_24_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_24_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_24_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_24_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_24_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_24_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_24_353 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_361 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_365 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_24_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_24_372 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_388 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_24_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_24_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_24_495 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_24_511 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_519 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_523 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_526 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_530 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_538 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_541 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_545 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_549 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_553 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_24_565 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_601 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_24_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_24_650 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_24_666 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_679 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_689 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_703 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_718 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_24_728 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_736 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_738 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_760 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_24_767 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_775 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_779 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_781 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_24_784 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_24_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_24_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_24_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_25_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_25_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_25_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_25_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_25_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_25_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_25_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_25_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_25_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_25_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_25_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_25_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_25_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_25_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_25_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_515 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_518 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_520 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_523 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_535 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_539 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_543 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_545 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_554 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_561 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_565 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_573 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_588 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_592 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_618 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_622 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_624 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_25_658 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_666 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_670 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_672 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_675 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_700 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_708 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_25_726 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_25_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_762 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_790 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_797 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_25_801 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_809 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_813 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_823 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_833 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_839 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_25_843 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_25_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_25_890 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_25_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_25_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_26_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_26_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_26_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_26_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_26_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_26_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_26_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_26_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_26_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_26_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_26_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_26_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_26_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_26_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_26_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_26_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_26_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_26_479 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_487 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_500 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_504 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_507 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_511 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_517 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_541 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_26_588 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_596 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_612 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_614 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_617 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_627 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_637 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_652 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_662 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_666 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_670 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_682 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_696 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_710 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_714 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_718 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_735 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_771 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_773 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_782 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_808 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_812 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_832 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_846 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_850 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_858 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_865 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_871 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_875 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_879 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_26_896 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_26_928 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_26_944 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_952 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_956 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_26_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_27_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_27_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_27_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_27_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_27_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_27_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_27_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_27_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_27_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_27_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_27_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_27_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_27_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_27_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_27_444 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_452 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_459 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_494 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_506 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_513 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_547 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_554 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_556 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_579 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_586 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_588 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_591 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_595 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_631 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_635 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_643 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_652 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_654 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_657 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_661 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_687 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_701 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_27_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_720 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_724 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_728 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_27_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_742 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_759 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_773 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_796 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_800 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_804 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_833 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_848 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_860 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_864 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_866 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_875 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_885 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_895 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_27_899 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_27_915 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_27_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_27_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_28_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_28_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_28_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_28_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_28_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_28_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_28_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_28_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_28_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_28_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_28_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_28_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_28_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_28_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_28_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_28_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_426 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_500 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_508 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_510 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_516 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_523 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_541 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_545 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_551 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_558 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_571 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_575 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_582 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_586 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_588 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_594 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_615 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_28_622 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_28_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_646 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_655 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_664 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_671 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_689 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_693 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_697 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_699 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_708 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_710 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_713 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_717 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_719 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_722 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_726 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_730 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_750 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_778 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_798 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_805 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_832 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_846 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_850 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_859 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_861 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_885 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_28_914 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_28_946 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_954 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_28_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_29_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_29_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_29_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_29_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_29_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_29_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_29_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_29_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_29_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_29_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_29_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_29_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_29_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_29_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_493 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_509 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_517 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_519 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_525 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_537 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_539 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_546 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_550 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_573 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_587 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_591 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_609 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_619 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_623 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_29_631 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_645 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_654 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_656 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_659 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_680 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_684 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_691 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_697 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_701 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_708 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_722 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_729 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_29_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_736 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_743 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_764 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_771 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_777 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_794 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_800 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_826 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_830 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_834 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_838 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_879 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_899 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_29_909 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_917 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_921 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_29_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_29_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_1016 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_2_1020 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_2_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_1091 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_2_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_2_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_1181 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_2_1188 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_1204 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_1208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_1239 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_1274 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_1278 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_2_1282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_2_1298 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_1306 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_1310 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_2_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_1390 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_1397 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_1449 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_1453 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_2_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_2_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_2_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_2_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_2_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_2_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_2_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_2_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_2_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_2_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_2_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_2_550 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_558 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_2_566 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_2_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_2_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_2_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_2_779 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_787 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_2_794 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_810 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_814 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_2_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_940 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_2_944 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_952 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_956 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_2_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_2_976 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_984 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_986 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_30_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_30_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_30_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_30_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_30_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_30_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_30_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_30_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_30_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_30_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_30_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_30_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_30_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_30_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_30_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_30_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_514 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_522 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_541 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_548 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_573 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_583 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_591 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_595 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_607 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_614 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_629 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_637 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_30_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_649 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_652 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_656 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_665 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_672 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_679 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_683 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_695 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_713 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_717 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_720 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_724 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_728 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_732 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_739 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_741 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_757 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_759 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_762 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_769 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_773 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_805 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_824 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_826 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_835 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_863 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_867 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_883 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_903 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_913 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_30_921 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_30_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_31_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_31_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_31_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_31_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_31_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_31_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_31_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_31_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_31_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_31_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_31_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_31_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_31_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_432 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_436 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_467 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_31_471 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_479 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_483 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_485 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_488 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_501 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_504 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_508 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_515 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_517 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_520 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_530 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_540 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_548 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_555 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_560 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_583 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_590 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_595 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_603 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_609 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_616 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_631 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_635 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_648 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_652 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_656 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_658 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_661 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_665 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_668 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_672 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_31_675 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_693 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_697 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_701 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_708 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_715 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_719 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_727 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_729 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_31_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_732 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_736 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_743 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_754 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_756 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_759 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_766 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_773 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_803 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_813 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_822 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_826 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_833 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_841 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_845 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_849 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_860 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_870 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_896 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_900 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_915 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_31_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_31_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_975 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_979 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_985 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_992 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_31_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_32_1014 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_1022 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_1026 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_32_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_32_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_32_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_32_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_32_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_32_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_32_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_32_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_32_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_32_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_32_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_32_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_32_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_32_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_32_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_32_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_32_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_479 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_483 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_490 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_494 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_498 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_502 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_509 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_513 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_561 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_568 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_582 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_586 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_594 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_601 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_611 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_618 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_620 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_629 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_637 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_648 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_652 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_654 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_657 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_666 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_683 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_32_687 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_695 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_713 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_32_717 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_727 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_731 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_735 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_742 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_750 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_754 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_758 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_762 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_766 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_770 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_774 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_778 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_803 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_813 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_821 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_825 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_829 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_836 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_840 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_856 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_860 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_869 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_884 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_895 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_32_921 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_990 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_994 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_32_998 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_33_1003 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_33_1013 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_33_1045 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_1061 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_33_1070 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_1134 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_33_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_33_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_33_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_1354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_1360 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_33_1364 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_33_1396 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_33_1412 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_33_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_33_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_33_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_33_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_33_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_33_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_33_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_33_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_33_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_33_444 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_452 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_502 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_530 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_532 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_541 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_548 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_573 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_575 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_589 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_599 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_607 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_609 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_623 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_630 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_637 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_650 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_654 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_660 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_664 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_668 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_683 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_687 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_689 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_706 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_715 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_725 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_33_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_733 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_33_741 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_749 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_755 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_763 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_765 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_795 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_799 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_808 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_812 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_816 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_826 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_830 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_834 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_836 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_867 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_871 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_880 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_894 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_904 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_916 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_33_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_941 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_943 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_973 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_983 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_991 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_999 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_1011 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_1015 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_34_1019 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_1027 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_34_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_1043 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_1073 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_1075 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_1078 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_34_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_1080 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_1083 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_34_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_34_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_34_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_34_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_34_1276 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_34_1292 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_1300 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_1304 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_1318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_34_1322 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_1330 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_1333 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_1337 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_1343 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_1347 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_1355 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_1359 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_1362 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_1366 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_1370 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_1374 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_1378 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_1382 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_34_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_34_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_34_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_34_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_34_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_34_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_34_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_34_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_34_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_34_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_34_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_34_479 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_487 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_490 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_503 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_513 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_523 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_530 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_547 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_551 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_555 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_573 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_577 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_584 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_609 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_619 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_633 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_647 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_655 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_662 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_679 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_683 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_686 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_693 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_708 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_717 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_34_721 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_729 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_741 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_34_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_763 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_766 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_770 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_774 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_782 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_788 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_796 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_800 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_814 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_827 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_831 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_835 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_839 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_843 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_861 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_863 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_872 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_34_878 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_905 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_938 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_942 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_946 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_949 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_35_1026 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_1034 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_1038 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_1042 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_1046 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_1050 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_1053 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_1055 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_1058 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_1070 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_1074 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_1077 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_1081 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_1085 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_1089 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_1093 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_1097 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_35_1103 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_35_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_35_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_35_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_1296 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_1300 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_1304 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_1316 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_1320 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_1326 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_1330 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_1333 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_1335 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_1338 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_1342 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_1354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_1358 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_1362 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_1366 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_1370 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_1373 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_1377 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_1381 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_1385 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_35_1389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_35_1405 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_1413 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_1417 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_35_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_35_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_35_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_35_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_35_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_35_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_35_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_35_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_35_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_436 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_440 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_442 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_445 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_476 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_480 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_494 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_503 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_507 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_511 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_519 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_523 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_526 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_530 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_532 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_535 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_539 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_545 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_552 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_575 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_589 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_604 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_608 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_617 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_629 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_631 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_655 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_659 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_675 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_679 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_683 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_685 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_688 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_695 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_708 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_715 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_721 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_727 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_35_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_35_731 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_739 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_743 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_35_746 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_762 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_766 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_770 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_774 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_790 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_800 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_808 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_817 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_848 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_856 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_869 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_871 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_874 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_908 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_916 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_920 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_35_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_943 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_951 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_959 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_969 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_979 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_983 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_1011 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_1018 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_1022 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_1026 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_1034 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_1038 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_1040 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_1043 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_1045 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_1048 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_1079 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_36_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_1083 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_1091 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_1104 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_1109 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_1113 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_36_1117 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_1125 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_36_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_36_1163 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_36_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_36_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_36_1276 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_1292 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_1296 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_1300 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_1304 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_1318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_1322 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_1326 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_1330 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_1334 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_1338 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_1342 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_1346 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_1350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_1354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_1358 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_1362 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_1366 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_1368 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_1371 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_1375 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_1389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_1393 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_1397 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_1401 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_1405 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_1407 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_1410 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_1414 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_36_1418 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_36_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_36_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_36_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_36_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_36_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_36_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_36_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_36_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_36_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_36_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_471 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_475 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_490 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_502 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_504 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_510 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_514 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_518 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_540 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_556 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_568 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_581 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_588 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_611 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_615 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_627 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_633 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_652 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_666 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_670 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_679 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_683 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_687 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_690 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_694 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_698 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_710 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_714 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_750 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_756 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_758 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_788 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_792 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_796 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_798 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_801 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_805 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_857 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_36_861 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_869 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_873 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_36_876 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_884 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_36_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_905 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_909 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_36_915 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_36_931 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_939 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_945 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_949 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_970 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_977 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_1005 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_1038 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_1042 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_1046 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_1050 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_1054 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_1062 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_1076 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_1078 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_1129 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_1134 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_37_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_37_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_1282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_1285 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_1287 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_1290 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_1294 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_1298 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_1300 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_1303 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_1307 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_1309 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_1316 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_1320 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_1324 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_1327 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_1333 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_1337 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_1341 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_1354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_1358 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_1362 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_1366 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_1372 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_1374 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_1377 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_1382 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_1390 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_1394 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_1398 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_1402 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_1406 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_1410 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_1414 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_1418 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_1425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_37_1429 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_37_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_37_1461 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_37_1477 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_1485 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_1489 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_37_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_37_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_37_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_37_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_37_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_37_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_334 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_338 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_341 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_345 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_347 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_366 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_37_370 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_37_402 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_37_418 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_37_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_37_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_481 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_505 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_509 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_517 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_538 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_541 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_545 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_552 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_579 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_595 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_613 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_617 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_624 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_671 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_675 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_679 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_682 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_692 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_719 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_725 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_37_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_754 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_758 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_769 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_834 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_838 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_844 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_37_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_37_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_902 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_906 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_908 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_911 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_915 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_919 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_955 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_959 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_963 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_970 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_974 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_978 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_980 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_983 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_987 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_991 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_1000 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_1002 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_1011 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_1015 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_1019 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_1023 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_1027 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_1034 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_1040 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_1050 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_38_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_1081 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_1091 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_1093 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_1098 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_1132 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_1136 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_38_1140 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_38_1156 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_1164 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_1168 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_38_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_38_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_1260 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_1263 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_1267 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_1271 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_1275 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_1279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_1285 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_1287 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_1290 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_1294 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_1298 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_1306 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_1310 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_1318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_1322 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_1324 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_1327 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_1358 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_1366 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_1370 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_1374 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_1378 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_1382 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_1389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_1393 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_1397 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_1401 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_1405 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_1409 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_1413 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_1417 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_1421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_1425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_1429 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_1433 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_1437 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_38_1441 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_1449 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_1453 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_38_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_38_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_38_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_38_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_38_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_245 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_38_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_38_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_298 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_38_301 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_38_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_339 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_341 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_38_363 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_38_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_38_379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_408 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_412 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_433 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_38_437 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_453 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_38_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_38_479 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_487 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_495 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_497 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_38_500 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_508 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_512 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_515 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_519 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_526 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_528 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_540 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_547 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_573 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_577 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_584 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_594 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_596 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_608 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_618 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_624 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_637 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_650 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_660 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_662 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_665 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_706 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_710 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_713 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_752 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_756 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_759 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_792 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_796 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_798 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_801 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_805 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_809 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_813 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_821 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_825 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_836 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_38_855 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_38_871 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_879 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_896 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_900 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_904 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_908 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_910 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_913 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_924 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_931 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_935 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_939 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_943 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_949 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_966 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_1003 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_1036 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_1040 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_1042 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_1051 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_1062 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_1076 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_1082 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_1084 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_1114 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_1118 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_1126 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_1130 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_1134 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_1140 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_39_1149 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_39_1181 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_39_1197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_1205 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_39_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_39_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_1249 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_1251 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_1254 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_1258 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_1261 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_1265 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_1269 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_1283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_1289 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_1293 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_1303 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_1311 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_1319 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_1321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_1328 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_1332 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_1342 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_1346 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_1358 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_1366 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_1370 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_1374 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_1387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_1391 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_1395 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_1399 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_1403 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_1407 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_1411 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_1425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_1429 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_1433 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_1437 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_39_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_1441 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_1445 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_1449 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_1453 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_39_1456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_1488 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_39_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_39_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_39_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_39_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_231 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_235 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_254 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_39_258 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_274 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_278 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_297 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_305 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_39_309 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_327 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_39_337 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_345 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_347 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_39_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_39_373 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_383 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_393 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_397 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_401 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_405 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_407 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_410 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_414 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_444 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_448 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_455 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_459 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_467 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_471 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_473 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_39_476 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_495 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_39_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_507 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_510 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_516 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_520 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_543 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_549 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_553 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_579 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_583 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_590 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_606 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_631 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_635 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_651 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_658 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_662 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_692 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_694 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_697 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_708 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_721 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_725 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_729 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_39_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_733 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_748 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_752 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_756 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_760 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_767 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_777 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_799 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_816 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_820 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_824 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_828 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_838 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_846 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_850 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_857 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_861 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_878 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_894 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_902 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_909 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_913 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_935 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_939 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_943 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_951 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_955 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_959 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_966 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_970 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_986 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_990 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_999 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_3_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_3_1083 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_3_1093 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_3_1125 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_1133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_3_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_3_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_1217 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_1227 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_1231 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_1233 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_1240 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_1251 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_1259 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_1267 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_1271 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_1275 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_3_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_3_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_3_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_1391 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_1395 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_3_1399 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_3_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_3_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_3_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_3_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_3_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_3_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_3_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_3_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_3_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_3_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_3_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_3_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_3_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_3_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_3_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_3_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_3_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_3_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_1003 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_1012 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_1016 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_1020 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_1036 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_1042 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_1046 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_1077 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_40_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_1081 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_1089 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_1153 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_1159 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_40_1163 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_40_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_40_1205 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_40_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_1229 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_1235 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_1239 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_1247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_1253 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_1257 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_1261 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_1265 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_1275 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_1281 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_1376 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_1380 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_1389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_1397 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_1401 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_1405 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_1423 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_1427 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_1431 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_1435 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_1439 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_1443 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_1447 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_1451 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_1460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_1464 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_1468 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_40_1474 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_40_1506 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_1522 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_40_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_40_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_40_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_195 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_40_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_201 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_211 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_40_214 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_222 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_226 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_229 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_231 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_234 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_246 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_257 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_261 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_264 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_268 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_274 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_40_278 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_294 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_296 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_40_299 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_40_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_329 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_331 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_334 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_40_358 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_40_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_40_374 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_382 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_386 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_408 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_418 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_424 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_427 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_431 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_438 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_440 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_443 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_453 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_474 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_478 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_482 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_485 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_493 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_500 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_502 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_508 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_516 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_522 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_529 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_537 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_543 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_547 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_571 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_573 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_584 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_592 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_599 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_612 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_614 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_617 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_648 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_650 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_653 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_670 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_679 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_731 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_735 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_40_750 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_758 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_760 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_763 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_767 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_778 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_784 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_40_788 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_796 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_805 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_821 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_825 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_838 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_846 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_852 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_856 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_860 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_864 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_868 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_885 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_892 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_896 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_900 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_906 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_913 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_920 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_924 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_963 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_973 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_981 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_995 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_999 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_1004 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_1013 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_1048 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_41_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_1063 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_1074 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_1133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_1140 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_1174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_41_1178 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_41_1194 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_41_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_121 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_1225 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_1227 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_123 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_1230 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_1240 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_1248 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_1250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_1257 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_41_126 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_1265 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_1311 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_1360 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_1368 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_1370 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_1400 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_1408 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_1416 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_1429 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_1437 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_41_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_1445 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_1449 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_1453 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_1461 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_1465 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_1469 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_1473 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_1477 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_1481 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_1485 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_1489 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_41_1496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_41_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_180 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_186 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_188 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_41_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_201 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_227 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_231 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_252 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_262 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_264 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_270 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_274 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_295 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_41_299 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_319 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_41_329 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_337 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_363 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_369 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_373 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_393 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_403 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_407 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_411 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_417 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_444 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_446 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_449 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_453 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_455 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_458 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_470 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_474 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_478 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_482 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_506 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_514 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_41_518 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_543 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_547 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_551 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_555 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_579 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_581 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_586 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_617 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_631 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_635 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_643 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_677 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_694 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_698 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_701 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_721 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_728 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_41_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_735 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_739 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_742 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_751 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_755 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_758 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_764 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_41_768 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_790 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_794 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_798 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_829 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_831 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_838 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_849 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_863 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_867 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_871 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_873 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_880 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_888 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_892 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_898 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_909 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_916 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_920 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_927 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_934 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_938 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_41_942 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_950 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_952 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_982 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_988 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_992 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_998 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_1010 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_1021 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_1025 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_1034 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_1036 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_42_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_1093 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_1111 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_1121 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_1125 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_1156 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_1176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_118 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_42_1180 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_42_1196 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_1204 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_42_1210 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_1218 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_122 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_1224 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_1228 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_1236 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_1238 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_1252 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_126 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_1283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_1291 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_1293 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_1302 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_1310 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_1322 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_1326 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_1328 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_1388 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_1418 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_1424 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_42_145 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_1460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_1464 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_1468 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_1472 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_1476 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_1480 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_1484 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_1488 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_1492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_1496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_1500 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_1504 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_42_1508 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_1524 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_42_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_153 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_156 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_42_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_162 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_186 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_197 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_42_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_201 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_217 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_231 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_239 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_254 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_260 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_268 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_275 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_292 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_298 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_302 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_306 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_42_310 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_42_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_339 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_341 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_344 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_358 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_360 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_363 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_367 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_42_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_374 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_378 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_380 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_388 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_395 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_399 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_403 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_405 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_408 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_412 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_42_415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_423 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_427 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_445 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_449 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_453 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_472 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_476 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_42_480 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_42_498 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_42_508 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_528 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_537 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_541 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_553 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_555 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_558 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_571 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_577 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_581 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_589 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_593 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_595 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_607 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_610 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_620 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_672 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_685 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_692 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_696 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_727 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_738 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_757 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_765 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_774 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_781 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_42_785 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_42_801 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_809 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_813 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_848 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_852 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_856 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_858 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_874 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_878 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_919 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_923 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_933 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_937 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_42_941 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_949 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_969 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_973 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_977 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_1038 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_1050 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_1062 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_1076 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_1078 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_1089 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_1093 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_110 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_1104 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_1116 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_1126 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_1130 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_1134 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_114 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_1140 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_1176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_118 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_1180 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_1184 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_1188 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_1196 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_1200 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_1239 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_1270 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_1274 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_1283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_1287 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_129 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_1296 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_1306 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_1314 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_1318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_1322 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_1331 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_1341 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_1360 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_1370 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_1372 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_1402 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_1406 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_1410 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_1424 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_1433 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_1464 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_1472 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_1476 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_1480 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_1484 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_1488 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_1500 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_1508 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_151 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_43_1512 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_43_1544 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_155 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_43_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_164 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_184 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_190 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_194 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_43_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_201 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_218 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_222 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_224 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_230 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_234 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_238 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_242 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_253 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_43_257 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_267 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_270 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_274 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_281 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_289 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_291 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_294 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_302 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_316 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_320 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_337 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_345 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_351 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_364 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_372 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_391 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_395 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_399 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_401 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_404 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_413 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_417 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_455 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_469 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_479 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_483 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_487 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_491 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_493 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_508 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_512 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_536 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_540 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_556 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_560 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_574 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_581 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_43_585 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_601 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_609 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_617 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_627 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_657 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_664 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_677 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_681 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_728 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_732 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_738 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_745 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_756 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_76 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_762 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_773 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_777 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_786 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_790 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_796 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_80 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_43_83 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_830 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_840 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_850 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_857 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_861 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_863 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_898 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_902 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_915 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_928 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_936 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_940 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_43_944 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_952 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_958 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_966 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_970 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_974 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_43_99 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_991 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_998 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_1011 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_1015 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_1019 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_1021 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_1061 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_1069 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_1077 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_1079 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_1086 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_1094 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_1098 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_1104 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_1111 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_1125 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_1139 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_1225 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_1227 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_1230 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_1234 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_125 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_1253 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_1263 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_1275 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_1305 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_1309 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_131 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_44_135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_1395 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_1405 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_1409 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_1421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_1452 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_1466 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_1474 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_1482 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_44_151 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_1523 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_44_1531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_44_1563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_1579 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_159 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_162 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_181 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_184 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_188 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_192 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_44_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_204 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_214 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_218 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_44_222 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_238 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_257 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_44_261 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_281 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_290 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_294 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_306 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_44_324 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_356 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_358 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_361 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_365 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_44_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_380 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_386 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_406 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_413 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_417 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_420 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_432 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_444 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_448 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_452 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_44_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_473 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_475 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_478 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_482 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_505 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_44_509 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_517 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_523 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_526 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_44_53 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_530 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_540 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_548 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_44_552 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_44_568 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_580 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_582 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_585 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_589 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_591 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_594 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_611 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_615 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_618 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_63 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_639 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_656 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_660 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_666 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_686 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_692 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_696 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_729 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_733 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_788 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_790 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_81 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_821 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_825 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_831 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_835 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_866 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_88 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_881 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_885 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_892 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_896 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_898 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_92 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_928 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_938 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_946 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_948 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_955 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_96 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_98 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_1029 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_1037 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_1049 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_1061 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_1076 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_1084 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_1092 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_111 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_1110 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_1114 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_1123 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_1133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_1141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_1143 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_1177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_1181 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_1185 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_1189 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_119 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_1193 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_1197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_1201 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_1205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_45_123 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_1239 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_1243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_1247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_1310 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_1318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_1326 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_1334 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_1346 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_1381 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_1389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_1397 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_1405 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_1413 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_1417 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_45_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_1473 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_1481 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_1489 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_1523 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_1527 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_45_1531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_45_1547 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_1555 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_1559 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_45_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_160 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_45_163 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_45_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_187 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_191 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_45_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_204 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_211 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_218 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_45_222 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_236 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_252 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_45_256 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_45_272 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_296 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_298 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_301 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_305 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_45_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_361 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_365 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_377 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_391 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_395 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_397 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_400 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_408 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_412 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_418 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_432 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_436 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_45_440 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_448 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_45_452 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_464 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_45_468 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_484 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_490 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_494 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_45_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_515 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_45_529 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_561 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_572 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_583 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_589 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_593 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_650 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_681 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_692 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_696 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_700 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_722 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_729 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_739 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_770 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_778 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_787 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_79 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_791 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_795 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_799 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_45_83 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_873 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_907 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_91 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_914 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_927 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_45_930 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_938 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_942 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_946 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_961 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_965 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_969 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_97 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_976 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_983 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_987 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_46_1002 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_1012 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_1018 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_1036 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_1038 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_1049 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_1059 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_1068 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_1077 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_46_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_1085 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_1091 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_1097 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_1105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_1109 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_1119 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_1129 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_1139 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_1149 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_1155 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_1161 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_1165 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_1169 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_1197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_1201 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_1205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_1216 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_1226 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_1236 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_46_124 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_1240 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_1295 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_1305 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_1309 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_132 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_1324 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_1357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_1367 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_1375 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_1393 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_1397 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_140 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_1409 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_1440 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_1448 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_1452 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_1470 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_1472 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_150 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_1502 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_1512 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_1520 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_1524 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_1531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_46_1535 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_46_1567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_1575 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_1579 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_161 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_165 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_169 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_46_182 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_46_198 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_46_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_216 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_230 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_46_234 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_242 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_246 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_254 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_256 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_262 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_46_266 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_288 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_296 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_300 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_304 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_46_308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_316 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_46_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_46_337 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_345 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_347 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_358 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_360 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_369 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_373 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_377 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_39 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_46_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_400 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_403 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_407 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_426 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_46_430 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_438 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_442 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_444 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_472 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_476 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_478 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_481 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_488 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_494 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_497 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_509 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_46_513 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_529 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_53 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_540 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_46_544 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_560 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_568 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_57 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_586 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_59 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_46_590 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_46_608 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_616 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_620 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_636 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_640 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_679 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_68 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_683 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_687 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_691 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_71 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_743 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_757 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_759 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_775 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_779 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_46_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_791 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_793 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_802 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_814 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_821 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_825 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_829 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_83 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_833 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_837 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_867 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_87 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_881 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_885 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_46_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_905 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_46_91 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_911 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_46_915 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_923 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_926 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_930 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_932 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_941 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_46_949 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_46_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_968 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_99 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_998 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_10 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_1007 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_1011 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_1013 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_1016 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_1020 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_1032 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_1051 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_1055 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_1075 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_1083 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_1089 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_1101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_1111 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_1115 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_1121 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_1125 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_113 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_1147 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_1155 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_1159 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_1163 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_47_117 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_1190 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_1204 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_1239 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_1247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_1259 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_1269 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_1287 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_1320 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_1328 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_1336 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_1354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_1369 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_1377 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_1384 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_14 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_1431 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_1462 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_1473 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_1477 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_1487 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_1495 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_150 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_1529 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_1533 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_1537 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_47_154 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_1541 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_47_1545 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_47_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_162 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_164 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_17 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_183 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_47_187 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_47_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_210 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_219 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_230 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_47_234 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_260 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_267 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_27 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_47_271 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_47_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_294 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_302 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_306 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_47_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_337 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_339 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_342 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_369 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_38 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_380 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_47_388 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_396 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_400 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_407 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_411 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_47_415 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_47_42 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_423 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_432 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_435 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_439 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_452 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_466 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_470 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_481 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_487 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_502 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_514 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_518 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_520 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_526 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_536 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_544 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_47_548 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_577 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_58 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_584 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_588 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_596 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_47_604 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_620 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_623 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_633 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_637 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_645 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_649 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_652 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_656 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_660 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_664 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_668 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_672 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_675 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_685 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_689 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_47_693 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_719 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_723 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_727 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_47_731 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_739 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_745 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_749 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_757 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_76 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_767 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_775 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_777 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_786 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_47_790 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_798 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_47_80 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_802 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_816 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_824 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_826 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_835 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_839 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_860 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_868 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_872 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_876 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_88 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_880 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_47_890 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_47_906 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_914 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_92 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_47_932 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_47_948 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_956 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_47_964 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_980 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_47_999 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_1000 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_1006 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_1014 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_1020 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_1049 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_1058 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_1062 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_1074 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_1082 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_1094 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_1098 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_1109 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_1113 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_1117 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_1121 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_1125 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_1134 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_48_114 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_1144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_1154 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_1197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_1228 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_1236 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_1240 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_1274 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_1282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_48_130 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_1324 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_1332 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_1336 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_1352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_1356 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_1380 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_1403 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_1407 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_1409 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_1439 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_1449 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_1453 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_1464 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_1472 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_1484 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_1492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_1523 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_48_153 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_1535 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_1539 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_1543 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_1547 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_48_1551 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_48_1567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_1575 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_1579 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_161 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_167 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_48_189 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_48_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_48_205 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_213 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_219 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_228 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_232 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_236 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_259 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_48_263 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_48_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_28 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_287 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_296 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_30 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_310 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_48_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_329 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_33 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_336 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_48_340 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_348 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_355 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_359 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_363 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_367 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_371 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_48_375 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_383 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_48_40 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_402 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_410 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_48_414 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_446 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_450 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_458 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_477 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_481 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_485 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_498 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_502 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_48_512 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_528 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_543 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_551 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_555 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_56 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_561 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_583 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_589 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_593 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_60 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_601 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_48_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_613 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_617 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_621 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_625 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_48_633 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_48_649 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_657 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_661 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_665 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_679 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_691 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_48_695 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_48_727 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_735 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_739 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_743 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_751 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_754 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_758 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_48_76 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_766 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_778 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_784 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_794 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_48_798 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_806 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_808 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_827 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_831 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_835 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_839 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_84 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_48_843 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_853 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_861 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_865 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_872 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_88 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_880 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_884 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_48_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_905 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_909 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_913 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_921 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_931 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_48_935 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_48_969 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_985 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_992 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_49_1003 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_1011 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_1015 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_1020 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_1032 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_1034 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_1041 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_1050 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_1059 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_1063 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_1074 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_1076 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_110 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_1105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_1113 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_1117 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_1119 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_1126 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_1134 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_114 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_1147 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_1155 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_1163 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_1167 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_49_118 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_1180 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_1194 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_1198 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_1212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_1216 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_1225 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_1229 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_1231 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_1252 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_1260 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_1271 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_1287 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_1295 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_1299 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_1332 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_49_134 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_1375 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_1377 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_1411 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_1432 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_1440 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_1471 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_1479 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_148 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_1487 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_1502 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_1506 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_1508 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_1559 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_156 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_49_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_164 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_169 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_180 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_49_184 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_194 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_49_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_200 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_204 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_22 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_49_223 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_239 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_24 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_252 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_49_256 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_49_272 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_297 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_307 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_31 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_49_315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_323 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_327 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_339 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_49_343 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_35 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_49_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_38 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_49_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_397 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_401 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_404 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_49_408 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_42 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_424 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_49_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_436 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_438 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_49_441 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_49_46 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_49_473 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_481 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_485 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_49_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_509 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_519 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_523 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_49_532 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_540 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_542 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_49_545 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_553 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_49_556 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_574 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_581 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_588 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_49_592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_608 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_612 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_619 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_49_62 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_636 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_49_645 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_677 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_686 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_694 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_49_698 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_706 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_717 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_721 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_725 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_751 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_49_755 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_763 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_765 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_768 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_49_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_790 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_794 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_49_80 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_824 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_828 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_841 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_845 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_849 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_88 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_90 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_905 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_49_909 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_917 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_921 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_929 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_93 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_933 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_952 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_956 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_49_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_97 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_49_976 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_984 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_988 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_990 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_4_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_1047 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_1049 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_1079 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_4_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_4_1083 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_4_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_4_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_4_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_4_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_4_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_4_1402 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_1410 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_1412 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_4_1442 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_4_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_4_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_4_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_4_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_4_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_4_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_4_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_4_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_4_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_4_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_4_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_4_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_4_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_4_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_4_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_4_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_897 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_901 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_4_932 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_4_948 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_956 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_4_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_50_1013 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_1021 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_1025 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_1036 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_1038 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_1045 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_1053 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_1066 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_1070 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_1084 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_1097 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_1112 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_1116 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_1120 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_1124 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_1126 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_1133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_1141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_1145 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_1161 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_1165 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_1169 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_117 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_1182 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_1184 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_1193 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_1201 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_1205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_50_121 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_1211 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_1218 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_1226 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_1230 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_1247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_1257 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_1261 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_1272 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_1276 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_1279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_1287 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_1295 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_1299 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_1325 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_1336 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_1345 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_1370 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_1378 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_1382 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_140 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_1411 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_1424 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_1451 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_1465 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_1469 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_147 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_1473 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_1482 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_1513 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_1523 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_1558 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_1562 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_50_1566 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_157 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_1574 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_1578 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_159 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_165 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_169 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_192 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_194 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_197 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_50_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_201 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_211 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_225 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_228 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_234 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_238 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_245 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_50_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_50_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_290 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_294 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_50_297 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_313 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_50_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_329 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_333 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_345 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_50_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_365 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_369 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_371 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_50_374 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_382 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_386 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_39 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_402 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_50_406 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_42 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_429 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_433 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_444 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_448 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_50_452 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_50_46 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_465 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_472 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_50_476 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_495 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_507 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_518 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_522 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_50_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_542 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_546 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_554 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_50_565 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_583 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_592 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_596 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_600 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_50_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_613 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_617 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_628 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_645 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_655 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_659 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_50_663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_671 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_50_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_684 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_688 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_50_692 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_700 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_707 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_715 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_725 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_729 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_733 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_735 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_741 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_50_758 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_50_78 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_50_792 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_50_808 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_825 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_829 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_833 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_837 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_839 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_869 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_871 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_50_878 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_50_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_50_905 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_913 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_917 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_50_929 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_94 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_50_945 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_50_963 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_50_979 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_98 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_50_997 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_51_1007 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_1023 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_1027 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_1029 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_1032 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_1036 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_1043 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_1055 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_1081 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_1089 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_1091 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_1103 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_1116 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_1120 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_1124 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_1128 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_1132 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_1145 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_1153 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_116 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_1160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_1164 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_1168 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_1172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_1176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_1180 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_1184 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_1188 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_1196 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_1200 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_1204 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_1212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_1216 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_122 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_1224 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_1232 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_126 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_1263 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_1271 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_1275 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_51_130 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_1331 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_1341 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_1353 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_1370 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_1397 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_1407 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_1411 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_1425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_1477 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_1481 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_1523 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_1531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_1539 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_1543 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_1547 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_1551 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_1555 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_1559 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_1567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_157 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_51_1571 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_1579 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_159 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_162 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_175 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_186 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_188 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_191 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_51_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_20 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_220 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_224 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_230 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_240 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_258 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_51_262 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_278 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_295 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_303 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_51_307 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_31 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_51_331 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_51_347 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_35 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_361 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_372 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_378 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_382 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_51_388 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_51_39 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_404 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_408 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_411 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_430 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_439 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_443 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_447 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_455 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_458 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_475 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_51_479 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_495 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_505 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_517 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_51_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_51_537 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_545 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_549 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_55 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_556 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_57 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_51_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_604 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_607 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_611 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_618 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_628 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_636 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_51_644 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_652 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_656 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_658 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_665 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_51_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_51_701 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_51_719 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_735 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_739 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_743 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_745 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_748 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_51_752 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_51_768 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_51_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_51_799 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_80 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_51_810 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_51_826 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_834 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_838 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_51_84 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_841 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_51_857 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_865 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_871 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_51_875 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_891 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_895 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_899 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_51_907 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_915 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_919 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_92 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_51_932 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_940 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_942 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_945 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_949 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_964 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_971 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_51_975 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_983 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_985 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_988 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_992 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_999 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_52_1003 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_52_1019 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_52_102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_1027 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_52_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_1041 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_1045 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_1049 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_52_1057 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_1066 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_1075 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_52_1081 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_1105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_1109 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_1113 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_1117 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_1121 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_1125 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_1129 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_1133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_1137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_1145 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_1149 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_52_115 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_52_1153 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_1159 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_1163 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_52_1167 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_1176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_1180 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_1184 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_52_1188 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_119 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_1196 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_1199 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_1203 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_1207 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_1211 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_1215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_1219 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_122 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_1231 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_124 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_1274 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_1282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_52_1290 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_1294 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_1301 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_1345 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_1352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_1360 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_1378 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_1382 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_52_1396 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_1429 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_52_1433 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_1437 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_1447 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_52_1451 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_1467 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_1475 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_52_1479 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_1483 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_1513 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_1531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_1535 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_1539 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_154 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_1543 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_1547 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_1551 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_1555 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_52_1559 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_52_1575 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_1579 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_52_168 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_175 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_182 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_52_186 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_194 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_197 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_52_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_201 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_219 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_22 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_52_223 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_52_239 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_245 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_52_262 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_52_294 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_308 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_52_312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_316 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_32 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_52_324 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_52_356 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_374 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_52_386 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_399 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_52_403 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_420 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_424 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_438 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_442 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_446 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_46 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_474 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_478 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_52_482 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_52_498 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_52_50 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_506 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_509 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_52_513 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_529 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_536 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_539 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_52_543 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_547 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_551 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_52_555 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_571 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_573 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_596 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_600 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_615 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_619 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_623 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_52_627 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_52_659 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_52_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_52_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_671 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_52_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_708 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_710 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_52_713 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_52_729 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_760 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_764 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_52_768 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_52_78 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_52_784 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_792 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_804 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_808 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_52_812 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_52_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_82 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_86 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_52_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_897 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_90 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_52_901 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_52_933 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_94 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_52_949 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_52_964 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_52_972 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_976 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_979 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_52_986 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_990 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_995 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_1012 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_1016 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_1018 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_1021 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_53_1029 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_1045 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_1049 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_1053 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_1057 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_1061 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_1077 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_1085 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_1093 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_1097 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_1101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_1105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_1109 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_1113 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_1117 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_112 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_1121 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_1125 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_1129 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_1133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_53_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_1154 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_1158 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_53_1162 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_1194 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_1198 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_120 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_1211 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_1214 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_1218 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_1222 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_1230 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_126 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_1261 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_1287 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_1295 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_1299 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_130 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_1329 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_1339 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_1347 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_1356 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_1387 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_1395 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_1399 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_140 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_1408 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_1418 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_1429 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_1433 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_1442 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_1452 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_1456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_1458 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_1467 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_1477 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_1481 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_150 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_1502 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_1512 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_1520 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_1524 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_1532 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_1536 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_154 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_1540 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_1544 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_1548 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_1552 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_1556 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_53_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_162 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_181 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_185 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_53_188 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_196 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_53_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_200 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_205 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_218 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_222 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_226 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_233 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_253 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_257 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_26 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_263 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_53_271 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_53_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_30 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_53_302 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_310 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_322 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_53_334 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_53_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_53_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_373 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_376 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_53_380 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_412 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_423 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_53_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_436 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_440 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_443 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_455 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_468 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_472 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_53_482 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_490 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_494 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_53_506 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_514 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_518 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_520 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_523 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_537 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_547 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_554 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_558 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_573 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_612 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_616 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_620 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_627 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_631 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_53_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_649 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_660 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_53_664 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_672 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_678 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_681 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_689 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_693 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_697 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_701 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_750 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_752 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_76 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_765 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_769 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_53_773 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_53_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_80 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_803 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_53_819 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_827 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_831 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_838 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_84 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_53_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_850 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_53_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_870 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_874 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_881 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_53_885 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_917 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_921 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_53_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_941 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_53_961 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_53_977 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_98 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_985 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_991 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_53_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_10 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_1002 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_54_1006 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_1022 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_1026 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_54_1036 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_1048 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_1050 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_1053 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_1057 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_1074 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_1078 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_1082 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_1086 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_1090 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_1094 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_1096 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_1109 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_1119 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_54_1123 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_1133 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_1141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_1145 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_1148 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_54_115 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_1156 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_54_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_1205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_1213 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_1217 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_1225 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_1229 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_123 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_1233 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_1250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_126 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_1260 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_1264 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_1295 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_1299 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_1303 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_1366 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_1376 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_1417 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_1421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_1467 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_1475 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_1479 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_1483 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_1513 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_1517 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_1531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_1535 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_1539 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_1543 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_1547 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_54_1551 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_54_1567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_157 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_1575 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_1579 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_159 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_162 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_166 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_186 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_192 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_54_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_200 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_204 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_207 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_211 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_214 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_218 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_222 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_225 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_229 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_253 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_26 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_263 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_267 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_54_271 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_30 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_303 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_305 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_316 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_324 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_328 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_331 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_54_343 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_351 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_353 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_54_360 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_54_376 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_388 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_54_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_400 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_406 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_414 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_418 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_54_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_441 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_445 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_54_466 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_48 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_482 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_500 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_54_508 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_52 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_54_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_54 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_541 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_547 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_557 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_54_561 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_569 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_57 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_573 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_577 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_585 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_595 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_61 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_615 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_619 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_54_623 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_54_639 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_64 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_647 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_649 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_652 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_668 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_672 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_54_679 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_687 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_54_691 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_701 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_707 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_711 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_54_715 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_731 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_735 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_739 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_743 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_749 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_752 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_756 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_54_760 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_54_792 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_80 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_54_808 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_54_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_54_850 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_866 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_87 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_870 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_874 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_892 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_54_896 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_54_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_920 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_924 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_931 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_935 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_54_945 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_95 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_974 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_54_978 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_994 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_55_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_55_1074 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_1084 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_1088 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_1091 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_55_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_1140 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_1149 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_1153 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_55_1161 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_1193 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_1197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_1199 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_1216 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_1220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_1224 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_1228 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_123 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_1236 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_1240 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_1251 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_1253 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_1256 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_126 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_1264 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_1268 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_1287 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_1295 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_1305 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_1325 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_1335 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_1346 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_1361 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_1392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_140 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_1400 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_1408 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_1416 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_1425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_1427 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_1488 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_150 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_1500 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_1508 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_1516 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_1520 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_1524 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_1532 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_1536 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_154 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_1540 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_1544 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_1548 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_55_1552 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_55_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_158 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_162 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_169 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_55_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_210 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_218 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_228 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_269 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_27 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_55_273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_281 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_55_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_294 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_298 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_55_306 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_55_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_55_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_373 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_55_380 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_396 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_400 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_402 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_405 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_417 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_55_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_55_464 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_55_480 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_488 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_55_510 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_55_526 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_53 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_538 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_542 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_549 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_55 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_556 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_55_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_578 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_58 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_582 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_584 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_587 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_55_591 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_62 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_55_623 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_631 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_633 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_636 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_645 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_647 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_55_650 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_682 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_689 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_693 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_695 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_715 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_55_719 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_727 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_741 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_745 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_55_748 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_55_764 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_793 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_55_797 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_55_813 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_82 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_821 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_824 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_828 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_846 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_850 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_55_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_86 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_870 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_874 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_878 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_888 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_55_892 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_90 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_55_908 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_916 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_920 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_55_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_94 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_946 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_950 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_954 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_956 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_959 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_55_963 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_97 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_55_979 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_987 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_991 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_55_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_56_1008 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_1016 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_1020 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_103 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_1035 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_56_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_1062 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_1065 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_1069 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_1077 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_56_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_56_1081 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_1097 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_1106 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_1108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_1111 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_56_1119 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_56_1151 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_116 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_1167 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_56_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_56_1189 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_1197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_1201 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_1204 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_1208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_1212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_1216 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_1220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_1228 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_1236 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_124 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_1240 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_1251 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_1255 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_1263 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_1267 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_1271 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_1290 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_1300 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_1304 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_1318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_1330 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_1334 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_1338 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_1345 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_1353 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_1361 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_1369 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_1373 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_1382 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_1393 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_1401 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_1409 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_1417 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_1421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_1428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_1436 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_1438 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_1445 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_145 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_1464 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_1468 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_1472 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_149 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_1523 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_153 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_1531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_1535 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_1539 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_1543 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_56_1547 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_157 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_1579 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_161 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_56_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_203 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_213 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_217 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_22 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_223 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_232 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_234 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_258 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_268 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_56_278 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_290 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_292 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_295 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_56_303 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_32 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_328 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_56_332 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_364 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_366 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_56_373 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_56_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_40 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_408 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_415 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_56_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_56_435 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_56_44 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_443 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_445 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_448 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_56_474 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_482 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_484 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_487 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_501 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_56_508 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_52 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_56_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_56_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_56_55 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_550 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_56_553 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_56_569 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_579 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_583 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_587 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_601 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_56_608 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_624 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_648 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_652 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_656 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_56_660 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_668 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_672 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_56_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_684 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_692 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_56_696 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_71 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_56_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_720 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_724 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_726 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_729 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_736 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_56_74 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_756 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_56_760 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_793 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_795 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_798 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_808 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_812 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_822 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_829 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_56_837 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_56_869 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_885 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_892 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_896 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_899 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_90 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_56_907 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_92 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_939 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_942 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_968 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_972 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_56_976 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_99 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_10 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_1005 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_57_1009 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_1041 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_57_1047 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_1055 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_106 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_1061 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_1074 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_1078 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_57_1091 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_110 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_1107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_1111 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_1121 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_57_1125 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_57_114 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_57_1145 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_57_1161 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_1169 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_1171 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_57_1174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_1182 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_57_1188 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_1213 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_1217 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_1229 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_124 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_1245 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_1253 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_1263 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_1267 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_1274 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_1287 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_1297 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_1301 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_1305 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_1313 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_1328 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_1332 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_1339 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_1358 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_1366 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_1370 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_1376 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_1380 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_1382 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_1396 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_1404 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_1412 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_1432 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_1463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_1467 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_147 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_1474 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_1482 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_1496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_1500 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_1504 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_1508 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_151 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_1512 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_1516 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_1520 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_1524 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_1532 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_1536 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_1540 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_1544 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_57_1548 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_1556 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_57_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_16 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_57_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_203 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_207 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_224 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_228 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_23 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_232 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_236 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_240 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_246 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_253 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_273 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_281 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_57_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_57_302 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_310 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_316 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_319 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_324 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_33 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_336 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_57_340 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_348 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_57_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_365 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_369 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_373 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_57_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_41 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_57_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_444 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_446 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_57_45 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_453 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_57_464 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_57_502 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_57_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_57_550 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_558 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_560 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_580 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_584 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_586 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_596 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_57_600 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_57_61 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_636 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_57_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_57_677 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_685 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_689 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_57_697 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_57_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_720 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_57_724 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_732 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_738 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_742 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_57_746 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_76 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_762 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_764 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_770 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_774 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_778 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_787 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_794 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_798 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_80 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_57_802 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_57_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_826 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_828 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_57_831 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_84 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_57_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_57_870 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_878 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_885 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_887 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_896 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_57_900 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_916 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_920 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_57_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_96 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_57_961 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_57_977 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_985 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_58_1003 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_58_1019 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_1027 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_58_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_1045 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_1053 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_1057 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_1071 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_1073 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_58_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_1082 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_1092 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_1096 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_1106 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_1114 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_58_1118 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_1150 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_1154 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_1160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_1164 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_1168 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_1180 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_1186 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_1217 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_1225 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_1235 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_124 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_1251 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_1259 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_1266 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_1270 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_1274 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_1281 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_1285 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_1289 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_1293 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_1303 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_1307 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_1311 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_1330 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_1340 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_1349 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_1353 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_1357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_1359 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_1368 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_1376 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_1437 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_1447 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_1451 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_1460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_1464 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_1468 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_1472 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_1474 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_1504 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_1508 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_1512 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_1516 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_1520 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_1524 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_1531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_1535 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_1539 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_1543 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_58_1547 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_155 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_157 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_1579 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_164 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_185 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_195 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_58_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_22 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_222 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_58_226 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_234 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_238 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_24 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_240 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_263 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_58_267 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_275 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_281 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_284 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_288 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_58_294 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_302 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_306 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_31 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_310 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_332 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_336 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_58_340 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_348 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_351 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_358 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_58_362 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_370 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_374 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_58_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_40 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_42 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_58_424 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_440 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_443 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_45 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_455 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_474 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_478 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_482 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_58_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_502 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_512 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_516 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_522 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_526 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_530 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_542 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_546 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_548 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_55 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_58_555 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_57 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_587 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_593 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_601 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_617 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_58_621 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_637 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_64 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_644 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_58_648 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_664 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_668 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_670 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_678 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_689 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_58_693 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_713 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_722 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_730 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_58_734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_74 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_742 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_58_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_779 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_785 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_58_788 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_58_804 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_812 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_58_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_58_82 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_58_834 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_844 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_850 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_58_858 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_876 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_883 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_58_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_90 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_58_921 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_58_937 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_945 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_948 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_952 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_956 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_58_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_97 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_976 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_58_980 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_988 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_992 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_999 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_10 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_1003 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_1007 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_59_1011 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_59_1027 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_1035 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_1047 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_1056 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_1069 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_1072 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_59_1076 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_1097 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_59_1101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_1119 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_1129 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_1133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_59_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_59_114 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_1204 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_1212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_1216 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_1220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_1224 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_1228 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_1238 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_1246 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_1250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_1254 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_1256 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_1262 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_1266 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_1270 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_1287 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_1295 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_59_130 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_1303 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_1311 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_1319 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_1323 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_1327 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_1331 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_1335 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_1339 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_1360 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_1370 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_1374 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_1380 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_1388 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_1396 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_14 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_1404 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_1408 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_1410 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_1417 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_1437 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_1468 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_1472 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_1482 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_1496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_151 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_1527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_1531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_1535 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_1539 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_1543 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_1547 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_1551 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_1555 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_1559 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_59_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_59_157 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_165 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_169 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_188 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_197 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_59_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_201 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_228 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_23 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_232 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_234 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_254 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_268 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_27 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_292 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_296 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_59_300 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_308 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_31 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_316 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_323 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_59_327 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_343 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_59_371 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_59_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_395 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_397 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_400 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_404 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_41 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_424 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_59_431 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_439 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_443 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_447 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_59_45 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_458 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_462 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_465 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_477 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_481 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_484 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_59_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_507 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_510 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_522 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_59_526 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_59_558 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_566 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_59_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_586 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_589 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_617 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_621 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_625 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_629 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_631 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_654 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_658 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_59_662 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_67 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_59_694 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_59_715 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_59_731 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_739 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_742 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_59_750 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_758 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_762 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_59_766 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_774 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_778 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_786 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_79 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_796 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_59_800 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_83 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_59_832 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_848 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_59_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_870 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_874 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_876 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_879 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_883 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_89 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_899 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_59_903 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_919 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_928 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_932 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_944 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_948 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_950 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_967 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_97 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_971 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_975 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_979 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_987 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_991 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_5_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_5_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_5_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_5_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_5_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_5_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_5_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_5_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_5_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_5_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_5_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_5_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_5_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_5_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_5_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_5_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_5_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_5_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_5_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_5_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_5_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_5_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_5_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_10 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_60_1006 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_1022 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_1026 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_103 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_60_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_1041 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_1045 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_60_1056 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_60_1088 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_1096 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_60_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_114 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_60_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_1189 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_60_1199 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_12 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_1207 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_1213 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_1217 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_122 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_1229 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_1256 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_60_126 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_1266 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_1270 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_1274 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_1276 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_1279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_1286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_1293 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_1301 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_1311 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_1321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_1328 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_1332 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_1336 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_134 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_1340 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_1352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_1356 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_1360 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_1364 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_1368 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_1372 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_1378 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_1382 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_1391 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_1395 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_1399 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_1403 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_1405 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_1435 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_1448 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_1452 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_1466 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_1468 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_1477 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_1503 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_1513 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_1517 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_1531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_1535 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_1539 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_1543 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_1547 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_1551 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_1555 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_1559 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_156 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_60_1563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_1579 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_160 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_60_164 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_60_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_187 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_189 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_192 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_60_196 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_60_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_204 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_21 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_223 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_234 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_238 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_240 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_262 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_269 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_291 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_299 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_60_303 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_31 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_325 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_60_329 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_337 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_60_341 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_60_361 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_377 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_388 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_60_395 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_60_40 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_403 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_407 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_410 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_417 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_60_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_60_453 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_60_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_473 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_485 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_497 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_501 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_508 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_510 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_60_513 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_529 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_537 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_541 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_548 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_552 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_60_556 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_572 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_576 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_60_579 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_58 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_60_595 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_609 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_60_613 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_60_645 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_60_661 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_60_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_60_692 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_700 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_711 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_718 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_722 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_60_726 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_60_74 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_742 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_751 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_753 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_762 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_769 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_773 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_775 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_782 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_791 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_60_795 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_834 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_838 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_60_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_850 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_856 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_866 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_60_870 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_60_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_90 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_921 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_928 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_60_932 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_94 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_940 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_944 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_946 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_60_949 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_96 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_60_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_60_976 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_984 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_988 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_99 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_990 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_997 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_61_1015 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_1023 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_1027 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_1029 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_1032 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_1036 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_61_1047 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_1063 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_61_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_1083 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_1086 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_1090 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_112 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_1121 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_61_1125 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_1140 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_1149 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_61_1153 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_1161 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_1165 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_1169 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_61_1181 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_61_1197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_1205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_122 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_1239 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_1249 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_1253 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_1260 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_1264 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_1268 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_1272 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_1276 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_1283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_1290 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_1298 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_1306 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_1313 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_1317 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_61_132 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_1327 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_1331 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_1335 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_1339 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_1343 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_1347 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_1353 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_1360 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_1364 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_1376 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_1380 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_1382 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_1391 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_1399 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_140 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_1407 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_1452 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_1456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_1460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_1462 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_1469 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_1477 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_1526 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_1530 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_1534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_1538 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_1542 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_1546 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_1550 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_1554 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_1558 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_61_1567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_1575 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_1579 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_61_181 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_197 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_61_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_20 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_61_204 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_222 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_226 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_23 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_230 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_234 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_242 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_246 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_252 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_256 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_258 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_61_269 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_281 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_288 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_297 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_301 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_304 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_316 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_327 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_33 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_337 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_343 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_347 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_61_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_61_373 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_61_396 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_61_41 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_61_412 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_420 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_424 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_432 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_435 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_447 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_61_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_459 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_470 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_474 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_478 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_49 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_490 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_511 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_515 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_517 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_520 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_530 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_540 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_61_544 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_55 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_560 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_577 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_581 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_61_585 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_61_601 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_615 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_619 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_621 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_624 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_636 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_61_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_67 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_688 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_692 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_61_696 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_704 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_708 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_61_715 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_61_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_75 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_755 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_759 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_761 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_764 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_61_768 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_61_78 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_61_786 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_824 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_61_832 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_848 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_61_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_890 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_894 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_898 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_61_908 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_916 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_920 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_61_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_94 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_959 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_962 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_966 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_61_978 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_98 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_61_999 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_10 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_1009 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_62_1013 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_1021 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_1025 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_1048 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_62_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_1070 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_1084 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_62_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_1187 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_1191 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_62_1195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_1203 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_1205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_1208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_1212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_1218 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_1226 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_1234 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_62_124 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_1256 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_1258 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_1288 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_1296 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_1298 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_1307 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_1311 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_132 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_1321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_1328 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_1332 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_1336 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_1346 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_1354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_1358 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_1362 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_1366 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_1374 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_1378 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_1382 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_1389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_1393 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_1397 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_14 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_1407 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_1409 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_1416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_1429 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_1442 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_1452 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_146 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_1487 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_1491 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_150 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_1522 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_1531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_1535 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_1539 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_154 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_1543 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_1547 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_1551 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_1555 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_1559 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_62_1563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_1579 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_162 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_183 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_185 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_188 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_62_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_21 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_219 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_236 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_240 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_281 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_285 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_289 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_296 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_62_300 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_316 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_62_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_329 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_343 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_62_355 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_62_371 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_382 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_40 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_401 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_62_405 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_62_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_429 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_435 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_439 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_44 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_455 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_459 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_470 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_62_474 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_48 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_62_506 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_52 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_62_522 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_530 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_62_537 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_62_553 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_575 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_585 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_62_589 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_59 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_601 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_607 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_610 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_622 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_640 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_643 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_647 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_668 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_672 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_62_679 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_62_695 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_703 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_713 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_717 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_729 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_62_733 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_741 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_62_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_76 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_62_763 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_771 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_773 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_62_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_62_792 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_800 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_804 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_806 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_62_821 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_83 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_837 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_841 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_848 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_62_852 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_87 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_898 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_906 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_62_91 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_910 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_914 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_62_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_926 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_930 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_937 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_62_941 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_62_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_62_976 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_984 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_99 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_990 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_994 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_63_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_1036 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_1040 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_1043 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_1051 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_1055 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_1059 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_106 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_1063 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_63_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_109 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_63_1103 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_63_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_1176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_63_118 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_1183 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_63_1187 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_1195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_1199 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_1216 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_1224 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_1231 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_1235 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_1243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_1256 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_126 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_1269 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_1287 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_1291 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_130 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_1322 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_1326 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_1328 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_1335 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_1381 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_1385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_1392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_1400 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_1408 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_1412 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_1429 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_1433 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_63_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_1463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_1467 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_1477 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_15 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_1502 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_1504 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_152 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_1534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_1538 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_1542 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_1546 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_1550 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_1554 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_1558 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_156 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_1567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_63_1571 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_1579 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_159 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_169 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_180 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_189 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_193 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_197 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_63_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_201 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_211 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_222 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_224 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_227 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_231 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_235 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_25 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_256 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_281 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_63_289 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_305 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_63_308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_32 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_340 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_342 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_63_345 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_353 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_63_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_36 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_378 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_382 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_63_393 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_40 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_63_409 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_417 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_430 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_436 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_438 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_44 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_444 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_63_448 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_63_464 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_472 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_63_478 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_48 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_494 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_63_502 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_510 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_63_513 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_52 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_545 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_549 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_56 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_561 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_565 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_63_584 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_63_616 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_63_626 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_63 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_63_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_67 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_63_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_681 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_685 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_689 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_697 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_63_701 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_63_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_746 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_749 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_753 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_766 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_774 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_778 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_63_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_799 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_80 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_803 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_805 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_63_808 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_63_824 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_834 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_838 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_848 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_63_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_86 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_63_870 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_878 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_90 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_911 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_63_915 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_63_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_94 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_941 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_945 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_63_949 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_63_961 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_98 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_63_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_100 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_64_1015 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_1023 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_1025 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_1038 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_1042 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_1050 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_1061 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_1065 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_1069 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_64_1073 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_64_1089 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_1111 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_64_1115 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_64_1137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_1145 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_1148 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_64_115 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_1150 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_64_1153 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_1161 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_1165 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_1167 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_1175 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_1205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_1213 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_1229 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_123 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_1236 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_1240 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_126 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_1274 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_128 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_1282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_1284 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_1296 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_1304 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_1322 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_1326 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_1356 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_1369 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_1377 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_1381 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_1389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_1393 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_1403 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_1416 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_1424 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_1428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_1432 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_1444 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_1460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_1464 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_1468 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_1472 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_1476 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_1480 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_1484 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_1488 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_1492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_1494 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_1503 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_1507 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_1511 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_1515 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_1519 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_1523 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_1579 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_158 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_162 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_64_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_64_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_230 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_242 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_254 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_261 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_278 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_28 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_64_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_294 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_298 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_306 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_313 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_32 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_64_324 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_356 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_359 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_363 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_367 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_64_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_383 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_64_395 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_403 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_407 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_411 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_64_423 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_431 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_435 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_64_438 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_476 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_478 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_481 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_487 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_498 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_509 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_515 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_519 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_64_523 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_53 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_64_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_56 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_566 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_578 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_586 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_64_590 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_60 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_64_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_637 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_643 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_64_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_692 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_64_725 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_741 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_64_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_76 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_64_779 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_787 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_789 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_792 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_796 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_806 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_813 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_82 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_64_821 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_64_855 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_64_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_89 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_64_905 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_913 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_917 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_919 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_926 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_93 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_934 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_938 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_941 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_945 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_96 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_64_967 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_64_999 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_10 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_1032 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_1036 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_1040 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_1048 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_1056 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_1070 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_1074 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_1078 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_65_1082 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_1114 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_1118 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_112 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_1126 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_1140 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_1146 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_1150 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_1152 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_116 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_65_1161 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_65_1177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_1185 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_1188 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_119 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_1196 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_1204 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_1216 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_1224 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_1226 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_123 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_125 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_1282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_1327 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_1340 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_1358 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_1366 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_1370 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_1374 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_1407 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_1417 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_1431 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_1483 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_1487 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_1503 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_1534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_1538 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_65_154 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_1542 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_1546 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_1550 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_1554 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_1558 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_65_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_162 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_188 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_65_192 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_65_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_211 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_218 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_222 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_228 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_232 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_236 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_246 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_252 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_256 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_26 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_264 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_274 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_278 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_290 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_294 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_298 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_302 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_320 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_65_324 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_332 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_65_338 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_65_365 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_65_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_391 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_397 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_401 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_41 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_414 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_418 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_65_435 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_443 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_447 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_449 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_65_45 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_452 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_466 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_65_470 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_65_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_494 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_502 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_506 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_514 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_518 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_65_529 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_65_545 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_553 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_65_556 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_65_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_65_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_61 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_610 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_618 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_65_622 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_63 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_65_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_657 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_661 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_65_674 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_65_690 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_698 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_721 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_65_725 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_741 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_745 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_749 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_753 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_765 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_65_769 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_777 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_65_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_65_799 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_810 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_814 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_823 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_65_827 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_84 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_843 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_65_864 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_65_896 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_904 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_908 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_91 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_65_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_920 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_65_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_93 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_65_941 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_949 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_951 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_954 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_96 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_961 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_65_965 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_981 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_983 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_988 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_992 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_65_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_1040 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_1054 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_1062 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_1069 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_1079 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_1083 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_1091 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_1097 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_110 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_66_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_117 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_1177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_1180 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_1184 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_1188 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_1231 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_1239 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_1247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_1255 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_1265 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_1269 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_129 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_1299 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_1306 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_1310 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_1318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_1322 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_133 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_1373 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_1377 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_1381 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_1389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_1391 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_1407 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_1421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_1423 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_1435 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_1448 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_145 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_1452 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_1468 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_1472 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_1476 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_1478 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_1485 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_66_149 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_1498 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_1511 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_1531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_1535 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_1539 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_1543 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_1547 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_1551 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_1555 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_66_1559 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_1575 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_1579 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_165 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_66_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_211 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_214 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_218 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_228 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_232 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_234 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_256 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_260 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_264 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_66_274 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_290 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_294 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_298 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_302 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_31 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_66_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_329 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_331 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_334 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_338 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_342 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_358 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_362 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_366 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_372 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_376 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_398 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_402 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_408 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_418 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_43 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_435 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_66_439 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_455 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_66_47 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_470 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_474 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_476 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_479 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_483 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_494 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_498 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_502 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_516 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_522 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_526 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_530 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_66_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_542 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_546 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_548 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_55 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_551 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_555 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_557 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_66_568 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_58 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_600 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_66_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_66_626 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_636 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_645 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_66_649 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_659 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_68 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_727 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_66_731 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_739 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_743 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_66_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_763 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_765 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_66_768 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_66_800 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_66_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_82 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_84 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_896 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_902 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_910 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_92 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_66_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_954 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_964 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_968 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_972 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_984 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_988 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_66_992 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_10 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_1002 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_1006 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_1015 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_1019 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_1023 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_1026 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_1030 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_1047 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_1051 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_1053 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_1062 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_1078 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_1082 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_1086 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_1090 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_1094 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_1096 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_1105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_1109 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_1113 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_1115 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_1118 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_67_1126 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_1134 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_67_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_114 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_67_1154 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_1162 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_118 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_1197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_1199 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_121 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_1211 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_1243 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_67_125 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_1255 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_1268 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_1276 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_1287 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_1295 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_1299 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_1303 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_1307 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_1311 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_1319 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_1323 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_1327 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_1337 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_1341 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_1345 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_1364 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_1372 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_1376 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_1380 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_1384 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_1388 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_14 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_1400 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_1406 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_1410 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_1412 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_1431 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_1435 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_1439 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_1452 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_1458 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_1462 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_1466 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_1470 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_1478 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_1501 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_151 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_1534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_1538 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_1542 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_1546 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_155 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_1550 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_67_1554 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_67_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_67_159 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_16 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_175 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_178 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_186 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_193 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_197 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_67_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_201 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_203 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_223 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_227 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_67_231 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_249 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_253 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_257 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_261 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_264 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_27 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_272 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_67_293 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_303 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_319 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_67_323 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_67_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_373 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_377 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_67_391 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_399 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_403 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_407 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_67_41 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_417 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_67_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_444 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_448 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_453 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_461 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_468 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_67_472 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_67_488 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_49 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_67_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_515 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_67_518 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_67_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_542 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_544 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_547 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_555 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_57 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_67_573 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_67_589 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_601 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_608 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_610 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_67_613 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_67_629 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_637 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_645 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_649 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_661 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_665 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_67_677 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_67_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_67_728 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_736 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_67_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_752 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_754 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_757 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_761 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_765 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_767 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_67_786 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_67_802 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_810 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_819 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_823 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_67_827 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_67_843 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_67_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_67_870 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_878 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_881 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_885 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_67_896 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_904 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_908 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_67_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_92 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_920 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_930 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_934 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_936 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_67_939 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_94 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_97 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_67_971 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_987 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_991 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_1000 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_1007 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_68_1011 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_1015 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_1020 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_1037 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_1046 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_1059 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_1069 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_1077 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_1084 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_1088 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_1092 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_68_1096 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_68_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_68_1118 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_68_1126 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_1130 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_1133 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_68_1141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_68_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_68_1165 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_1169 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_68_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_68_1181 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_68_119 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_1235 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_68_129 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_1296 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_1300 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_1304 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_68_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_1325 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_1329 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_1333 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_1335 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_1347 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_1361 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_1365 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_1369 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_68_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_1377 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_1381 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_1397 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_1401 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_1403 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_1433 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_1441 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_1443 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_1464 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_1468 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_1472 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_1476 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_148 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_1480 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_1484 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_1497 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_1507 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_1517 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_68_152 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_1531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_1535 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_1539 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_1543 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_1547 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_68_1551 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_68_1567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_68_1575 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_1579 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_68_168 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_68_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_68_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_183 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_185 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_68_188 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_68_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_68_204 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_68_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_225 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_68_229 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_68_237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_253 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_68_257 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_26 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_68_271 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_68_287 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_29 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_68_295 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_310 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_68_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_33 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_68_337 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_68_345 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_355 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_365 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_68_369 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_68_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_68_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_68_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_41 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_43 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_68_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_46 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_469 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_473 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_68_477 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_50 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_68_509 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_68_517 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_68_528 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_68_537 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_68_54 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_553 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_68_557 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_68_589 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_68_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_60 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_601 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_68_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_611 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_615 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_68_625 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_64 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_68_657 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_68_665 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_682 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_68_686 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_68_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_710 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_717 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_721 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_68_725 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_733 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_736 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_74 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_763 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_775 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_779 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_68_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_68_799 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_68_80 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_803 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_813 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_821 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_68_825 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_68_857 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_86 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_68_873 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_881 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_885 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_68_892 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_68_898 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_68_90 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_68_908 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_914 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_926 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_930 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_934 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_938 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_94 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_940 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_949 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_68_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_68_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_68_968 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_97 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_974 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_68_982 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_998 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_1012 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_1016 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_1019 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_1023 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_1033 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_1043 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_1051 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_1076 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_1083 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_1091 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_69_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_1115 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_1125 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_1129 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_1133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_69_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_69_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_1180 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_1188 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_1194 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_1198 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_1216 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_1224 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_1232 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_1240 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_1248 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_1252 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_1264 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_1268 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_1270 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_1295 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_1299 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_1303 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_1310 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_1341 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_1345 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_1360 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_1362 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_1373 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_1391 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_1395 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_1406 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_1414 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_1418 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_1425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_1435 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_1445 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_1453 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_1461 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_1465 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_1469 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_69_147 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_1473 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_1477 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_1496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_1498 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_1532 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_1536 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_1540 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_69_1544 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_69_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_69_163 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_175 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_178 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_191 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_195 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_69_199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_69_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_207 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_217 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_272 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_69_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_69_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_36 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_361 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_367 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_371 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_69_375 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_383 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_69_396 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_412 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_414 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_423 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_69_431 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_69_447 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_455 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_459 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_461 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_69_464 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_472 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_69_478 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_48 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_69_488 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_50 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_501 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_69_504 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_69_520 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_528 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_53 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_532 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_536 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_546 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_550 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_69_554 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_566 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_69_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_586 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_589 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_599 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_603 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_69_607 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_63 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_644 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_69_648 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_69_664 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_67 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_672 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_674 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_677 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_685 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_69_689 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_718 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_722 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_69_726 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_69_742 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_750 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_754 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_757 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_76 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_769 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_773 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_69_794 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_810 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_814 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_816 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_69_819 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_69_835 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_843 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_856 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_86 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_862 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_69_866 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_874 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_883 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_891 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_895 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_897 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_906 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_916 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_92 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_920 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_928 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_932 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_936 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_938 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_69_941 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_96 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_69_973 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_69_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_6_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_6_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_6_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_6_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_6_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_6_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_6_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_6_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_6_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_6_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_6_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_6_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_6_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_6_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_6_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_6_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_6_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_6_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_6_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_6_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_6_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_6_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_6_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_6_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_70_1000 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_1016 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_1020 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_1042 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_1055 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_1057 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_1068 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_1076 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_1080 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_1084 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_1088 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_70_1092 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_1104 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_70_1107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_70_1139 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_114 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_1149 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_1153 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_70_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_1189 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_1193 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_1196 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_1204 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_1210 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_1247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_1255 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_1263 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_1267 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_1271 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_1284 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_1288 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_1292 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_1296 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_1300 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_1304 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_1318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_1322 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_1324 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_1335 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_1347 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_1355 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_1359 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_1366 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_1370 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_1374 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_1378 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_1382 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_1393 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_1401 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_1409 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_1413 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_1417 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_1421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_1425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_1433 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_1447 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_145 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_1451 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_1464 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_1468 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_1472 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_1476 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_1480 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_1484 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_1488 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_1492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_1504 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_1508 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_1512 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_1516 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_1520 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_1524 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_1531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_70_1535 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_70_1567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_1575 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_1579 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_182 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_70_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_22 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_236 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_240 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_70_253 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_26 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_327 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_70_331 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_365 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_372 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_70_376 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_388 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_70_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_40 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_408 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_412 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_70_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_44 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_70_441 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_449 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_453 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_476 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_480 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_490 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_495 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_502 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_509 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_511 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_518 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_70_522 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_530 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_70_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_70_550 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_558 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_70_566 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_574 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_578 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_70_586 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_609 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_61 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_70_616 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_624 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_627 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_631 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_640 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_650 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_70_654 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_680 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_683 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_687 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_691 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_697 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_706 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_716 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_724 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_70_728 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_70_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_763 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_767 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_70_771 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_80 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_70_803 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_829 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_70_833 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_84 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_70_865 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_88 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_881 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_885 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_70_893 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_90 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_901 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_907 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_924 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_93 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_70_931 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_70_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_969 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_97 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_973 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_977 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_983 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_992 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_10 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_100 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_1030 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_1034 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_1038 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_1041 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_1045 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_1049 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_1059 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_1063 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_1070 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_1074 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_1078 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_71_1082 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_1090 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_1094 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_1105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_1113 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_71_1117 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_1133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_71_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_115 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_71_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_1178 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_1182 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_1186 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_119 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_1194 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_1198 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_122 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_1239 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_1243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_1247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_1251 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_1265 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_1283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_1291 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_1295 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_1299 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_1316 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_1320 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_1324 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_1328 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_1332 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_1336 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_1340 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_1358 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_1366 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_1370 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_1374 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_1381 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_1385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_1387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_1396 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_1410 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_1414 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_1418 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_1425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_1429 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_1435 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_1458 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_1462 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_1466 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_71_147 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_1470 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_1474 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_1478 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_1482 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_1502 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_1504 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_1534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_1538 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_71_1542 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_155 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_1558 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_71_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_159 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_161 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_164 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_71_180 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_71_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_20 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_71_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_231 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_235 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_71_238 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_71_270 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_278 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_28 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_71_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_302 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_71_308 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_316 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_71_32 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_325 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_331 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_342 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_71_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_71_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_71_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_40 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_71_405 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_71_415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_423 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_71_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_71_462 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_48 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_494 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_501 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_71_504 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_52 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_71_520 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_528 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_530 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_71_533 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_549 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_553 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_56 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_573 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_71_577 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_71_593 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_60 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_601 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_603 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_606 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_71_614 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_630 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_653 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_71_657 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_671 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_681 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_688 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_690 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_699 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_703 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_707 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_714 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_717 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_724 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_71_755 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_765 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_769 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_773 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_777 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_71_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_80 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_84 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_86 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_866 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_870 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_71_874 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_89 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_906 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_920 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_928 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_93 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_932 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_934 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_937 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_71_945 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_71_977 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_71_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_1040 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_1048 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_1056 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_1068 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_72_1072 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_72_1088 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_1096 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_1104 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_1107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_72_1119 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_112 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_72_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_1143 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_1147 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_1151 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_1155 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_72_1176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_1194 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_122 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_1224 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_1232 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_1236 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_1238 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_1248 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_126 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_1267 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_1279 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_72_130 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_1310 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_1326 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_1330 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_1334 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_1338 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_1346 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_1360 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_1368 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_1376 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_1380 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_1393 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_1401 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_1409 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_72_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_1413 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_1417 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_1421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_1425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_1429 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_1433 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_1446 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_1468 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_1472 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_1476 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_1480 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_1484 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_1496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_1509 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_1519 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_1523 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_1531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_1535 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_1539 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_1543 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_72_1547 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_1579 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_72_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_72_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_72_211 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_72_227 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_235 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_72_238 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_246 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_72_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_266 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_269 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_287 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_293 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_297 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_304 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_72_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_72_353 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_361 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_365 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_368 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_72_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_375 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_72_379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_72_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_400 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_404 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_413 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_418 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_426 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_434 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_72_438 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_458 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_471 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_72_475 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_72_507 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_515 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_518 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_537 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_72_541 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_560 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_575 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_72_581 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_601 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_72_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_680 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_684 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_696 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_700 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_731 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_741 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_75 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_753 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_757 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_769 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_72_787 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_72_79 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_795 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_799 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_72_803 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_822 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_825 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_72_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_885 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_72_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_72_921 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_72_937 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_945 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_95 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_951 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_955 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_72_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_72_976 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_984 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_988 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_99 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_990 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_100 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_1003 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_73_1007 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_1011 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_1015 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_1027 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_73_1035 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_73_1051 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_1055 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_73_1058 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_1062 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_73_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_109 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_73_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_73_1109 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_73_1125 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_113 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_1133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_73_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_73_1146 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_1150 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_73_1153 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_73_117 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_73_1185 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_73_1201 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_1205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_1239 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_73_1243 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_73_125 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_1258 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_1271 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_1275 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_1283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_1287 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_1289 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_129 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_1301 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_73_1305 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_1309 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_1322 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_1326 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_1330 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_1334 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_1338 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_1342 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_1346 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_1359 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_1367 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_1375 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_1387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_1389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_1400 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_1408 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_73_1416 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_73_1425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_1440 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_1453 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_1461 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_1465 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_1469 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_73_147 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_1473 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_1477 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_1523 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_1554 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_73_1558 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_73_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_163 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_167 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_73_175 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_73_183 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_187 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_73_190 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_73_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_73_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_210 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_73_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_219 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_224 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_73_236 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_242 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_73_246 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_278 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_297 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_301 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_303 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_73_306 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_73_338 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_73_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_73_370 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_73_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_403 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_405 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_414 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_73_418 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_73_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_436 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_73_439 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_455 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_464 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_73_468 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_476 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_479 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_488 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_73_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_73_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_73_539 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_543 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_545 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_548 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_552 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_73_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_566 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_73_579 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_585 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_73_589 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_73_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_613 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_615 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_73_624 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_73_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_636 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_73_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_645 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_647 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_654 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_658 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_73_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_73_662 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_672 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_679 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_73_683 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_73_699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_707 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_719 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_73_723 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_739 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_73_743 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_76 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_73_788 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_796 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_799 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_73_80 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_803 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_813 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_73_817 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_73_825 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_829 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_831 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_834 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_844 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_73_848 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_73_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_73_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_73_894 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_898 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_904 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_908 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_73_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_920 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_73_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_73_933 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_937 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_940 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_949 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_73_96 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_961 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_73_965 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_73_981 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_1015 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_1019 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_1023 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_1027 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_74_1043 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_1059 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_1062 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_1072 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_1076 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_74_1080 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_1096 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_74_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_74_1134 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_1142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_1145 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_1149 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_74_1176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_120 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_1208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_124 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_1259 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_1269 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_74_128 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_1281 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_1285 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_1289 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_1293 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_1300 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_1302 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_1309 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_1326 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_1330 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_1334 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_1350 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_1362 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_1372 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_1376 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_1393 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_1395 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_1407 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_1411 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_1423 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_1468 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_1472 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_1476 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_1478 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_1485 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_1489 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_1501 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_1509 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_1513 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_1517 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_1531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_1535 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_74_1539 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_74_1571 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_1579 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_74_160 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_188 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_194 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_74_198 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_74_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_74_214 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_22 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_222 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_226 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_24 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_74_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_74_27 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_74_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_290 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_294 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_296 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_74_299 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_307 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_74_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_74_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_353 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_359 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_74_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_370 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_374 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_74_378 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_74_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_400 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_404 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_407 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_415 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_74_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_437 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_445 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_449 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_45 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_453 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_74_471 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_49 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_74_503 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_511 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_515 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_517 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_523 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_53 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_74_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_57 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_74_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_74_637 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_645 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_74_651 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_671 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_74_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_799 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_80 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_803 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_813 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_74_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_74_84 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_900 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_904 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_74_908 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_92 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_74_940 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_956 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_96 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_74_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_976 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_978 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_981 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_10 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_100 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_75_1076 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_109 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_1108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_1110 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_1113 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_1117 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_112 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_75_1126 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_1134 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_75_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_75_116 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_75_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_1186 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_1196 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_1200 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_1204 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_75_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_1217 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_1219 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_1249 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_1264 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_1272 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_1276 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_1283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_1287 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_1291 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_1293 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_1296 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_75_132 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_1327 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_1335 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_1343 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_1347 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_1358 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_1362 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_1366 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_1396 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_1398 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_14 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_140 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_1407 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_1425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_1438 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_75_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_1469 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_1473 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_1477 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_1479 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_1505 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_75_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_16 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_168 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_178 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_182 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_190 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_194 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_75_198 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_75_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_210 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_75_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_231 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_235 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_75_239 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_249 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_25 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_252 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_256 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_263 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_75_267 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_75_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_302 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_306 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_31 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_310 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_325 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_329 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_75_333 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_75_35 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_353 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_75_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_75_373 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_75_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_75_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_444 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_452 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_458 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_75_466 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_75_482 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_490 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_494 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_75_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_535 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_539 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_75_543 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_551 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_75_555 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_75_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_578 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_582 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_584 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_587 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_594 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_75_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_606 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_610 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_617 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_75_621 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_629 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_633 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_635 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_647 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_657 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_75_661 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_67 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_677 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_681 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_685 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_75_694 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_722 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_75_726 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_742 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_746 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_749 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_753 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_757 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_75_76 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_763 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_775 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_779 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_75_786 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_75_802 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_810 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_75_820 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_75_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_75_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_75_902 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_75_92 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_920 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_75_928 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_75_944 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_952 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_75_964 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_75_980 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_988 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_992 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_75_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_76_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_1027 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_76_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_76_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_76_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_76_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_1134 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_76_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_1175 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_76_1178 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_76_1194 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_1198 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_1200 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_1203 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_76_1211 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_1219 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_76_1226 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_1230 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_1233 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_76_1247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_1251 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_1263 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_1271 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_1279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_1283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_1287 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_1291 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_1295 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_1297 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_76_1309 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_1366 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_76_1398 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_1408 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_1416 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_1420 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_76_1451 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_1460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_1464 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_1468 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_1472 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_1476 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_1484 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_1488 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_76_1519 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_1523 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_76_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_76_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_76_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_76_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_76_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_76_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_254 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_266 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_76_270 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_76_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_290 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_294 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_76_308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_76_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_76_329 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_333 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_335 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_338 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_342 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_356 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_360 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_76_364 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_368 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_76_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_371 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_76_379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_76_403 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_76_435 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_76_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_458 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_466 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_470 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_76_480 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_76_498 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_506 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_513 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_517 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_536 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_539 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_543 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_553 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_76_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_599 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_611 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_76_615 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_76_647 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_76_663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_671 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_76_683 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_699 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_76_706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_76_738 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_742 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_76_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_753 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_765 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_76_769 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_76_801 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_76_809 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_813 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_76_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_76_834 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_845 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_76_856 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_864 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_76_868 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_884 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_896 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_76_900 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_904 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_907 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_76_911 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_921 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_76_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_76_941 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_949 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_956 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_76_963 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_77_1004 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_1008 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_77_1012 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_1020 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_77_1032 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_77_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_77_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_77_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_1151 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_77_1155 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_1165 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_77_1169 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_1176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_1185 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_77_1189 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_119 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_1205 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_77_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_1225 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_123 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_77_127 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_1310 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_77_1314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_1318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_77_135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_1381 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_1389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_1397 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_1399 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_1406 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_1431 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_1433 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_1442 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_1452 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_1456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_1460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_1464 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_1468 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_77_1472 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_1482 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_1496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_1500 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_1504 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_1508 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_1512 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_77_1516 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_77_1548 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_77_1556 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_77_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_175 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_77_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_77_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_183 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_185 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_190 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_77_194 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_198 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_77_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_201 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_77_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_77_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_223 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_226 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_236 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_240 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_77_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_77_26 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_77_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_77_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_30 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_302 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_77_305 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_77_313 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_32 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_77_320 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_77_336 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_342 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_77_360 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_77_376 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_77_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_39 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_423 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_77_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_77_43 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_77_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_77_468 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_472 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_476 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_502 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_77_506 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_77_522 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_530 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_77_533 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_77_541 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_545 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_547 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_554 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_77_558 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_566 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_77_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_77_586 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_77_59 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_607 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_616 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_77_620 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_636 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_77_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_77_67 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_77_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_77_689 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_697 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_77_701 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_707 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_77_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_77_718 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_728 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_77_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_77_736 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_77_768 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_77_790 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_77_822 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_77_838 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_77_846 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_850 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_77_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_858 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_77_861 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_875 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_77_879 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_77_887 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_893 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_897 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_907 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_77_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_77_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_77_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_1000 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_1004 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_78_1008 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_1022 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_1026 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_1037 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_78_1041 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_78_1049 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_1053 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_1055 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_1058 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_1062 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_1074 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_1078 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_78_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_78_1082 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_78_1090 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_1094 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_1096 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_78_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_78_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_78_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_78_1205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_1213 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_1217 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_1225 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_1233 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_78_1247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_1251 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_1263 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_1267 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_78_1271 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_1275 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_78_1305 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_1309 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_1327 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_1340 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_1352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_1393 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_1397 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_78_140 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_1401 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_1432 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_1445 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_1449 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_1453 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_78_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_148 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_1494 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_1498 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_150 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_78_1502 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_78_1518 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_78_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_78_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_78_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_161 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_78_165 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_78_173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_78_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_78_195 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_78_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_220 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_78_224 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_78_240 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_78_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_78_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_290 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_293 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_303 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_307 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_309 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_324 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_78_328 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_78_344 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_78_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_78_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_370 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_377 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_78_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_78_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_78_408 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_414 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_423 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_426 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_436 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_440 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_78_444 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_78_452 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_472 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_78_476 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_484 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_78_487 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_78_503 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_78_511 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_78_517 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_78_525 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_529 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_78_53 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_78_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_552 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_568 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_78_572 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_78_594 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_609 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_61 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_611 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_621 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_625 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_78_629 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_63 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_78_661 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_78_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_78_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_680 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_78_684 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_690 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_698 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_700 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_716 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_723 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_78_727 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_735 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_78_754 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_78_786 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_78_80 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_78_802 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_806 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_808 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_813 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_78_821 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_829 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_831 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_834 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_846 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_850 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_852 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_859 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_78_867 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_78_883 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_78_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_905 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_78_909 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_78_941 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_78_96 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_78_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_964 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_968 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_988 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_992 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_78_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_79_10 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_79_1004 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_1008 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_1011 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_1018 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_79_1022 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_1026 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_79_1030 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_79_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_1062 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_1074 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_79_1078 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_1086 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_1088 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_1091 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_79_1111 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_79_1127 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_79_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_79_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_118 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_79_1186 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_1196 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_79_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_122 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_1254 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_79_1258 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_79_126 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_1262 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_1264 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_1267 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_79_1271 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_79_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_1290 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_1298 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_1300 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_1303 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_1307 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_1323 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_1331 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_1335 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_1363 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_1394 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_1398 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_14 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_1402 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_1406 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_146 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_1473 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_1477 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_1481 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_1485 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_1489 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_79_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_1497 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_1501 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_79_1553 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_79_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_157 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_79_161 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_79_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_79_187 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_79_195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_79_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_20 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_211 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_218 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_79_222 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_79_238 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_24 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_248 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_79_252 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_260 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_262 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_79_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_79_28 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_281 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_79_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_79_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_79_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_38 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_79_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_393 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_395 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_401 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_405 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_79_409 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_79_42 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_79_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_79_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_79_468 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_472 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_474 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_79_483 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_79_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_493 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_502 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_79_515 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_79_525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_79_541 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_79_549 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_553 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_556 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_79_564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_79_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_574 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_79_58 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_79_582 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_79_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_611 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_619 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_79_623 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_631 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_79_645 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_79_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_79_661 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_671 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_674 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_682 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_79_693 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_697 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_700 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_79_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_79_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_79_728 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_79_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_732 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_734 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_79_764 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_794 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_804 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_79_808 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_79_840 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_79_848 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_79_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_79_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_79_929 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_79_937 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_941 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_945 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_79_949 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_79_981 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_79_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_79_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_7_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_7_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_7_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_7_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_7_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_7_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_7_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_7_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_7_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_7_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_7_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_7_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_7_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_7_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_7_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_7_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_7_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_7_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_7_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_7_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_7_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_7_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_7_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_80_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_80_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_80_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_80_1063 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_1071 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_1073 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_80_1076 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_80_1092 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_80_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_1110 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_1112 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_1115 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_80_1125 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_115 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_80_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_80_1165 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_1169 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_80_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_80_1181 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_1185 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_1187 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_80_119 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_1190 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_1194 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_1211 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_80_1215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_1225 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_1228 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_1236 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_1238 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_1251 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_1255 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_1259 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_80_1263 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_1269 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_1281 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_1289 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_1293 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_1295 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_80_1298 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_1304 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_1322 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_1330 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_1332 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_1339 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_1347 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_1355 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_1357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_1369 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_1382 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_1393 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_1401 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_1405 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_1413 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_1423 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_1460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_1462 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_80_1492 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_80_151 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_1524 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_80_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_80_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_80_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_80_159 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_169 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_80_173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_80_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_189 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_80_193 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_80_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_80_225 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_80_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_245 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_80_263 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_269 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_80_273 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_80_289 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_293 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_295 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_301 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_80_305 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_80_313 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_80_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_334 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_80_338 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_80_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_80_370 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_378 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_380 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_80_383 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_80_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_408 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_418 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_80_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_80_43 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_80_438 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_444 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_466 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_80_470 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_80_478 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_482 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_80_485 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_501 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_504 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_512 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_519 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_80_523 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_80_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_544 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_548 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_555 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_571 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_80_575 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_583 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_592 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_80_596 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_80_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_80_615 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_80_631 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_635 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_643 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_80_651 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_80_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_671 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_80_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_682 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_684 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_690 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_80_694 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_726 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_729 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_733 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_80_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_80_75 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_757 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_80_765 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_80_797 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_813 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_80_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_80_826 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_832 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_840 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_80_844 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_85 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_80_876 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_927 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_80_93 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_80_943 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_956 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_80_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_81_100 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_1012 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_1014 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_1021 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_81_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_81_1047 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_81_1055 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_1059 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_1061 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_1074 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_81_1082 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_110 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_1114 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_1117 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_1121 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_81_1129 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_1133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_81_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_1148 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_1162 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_81_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_81_1198 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_81_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_81_1225 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_1231 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_1239 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_81_124 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_1247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_1249 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_1256 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_1260 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_1296 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_1304 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_1339 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_1347 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_140 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_81_1402 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_1406 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_1412 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_1430 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_1432 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_81_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_1444 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_1464 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_1468 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_81_1472 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_1488 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_81_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_81_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_81_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_160 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_81_164 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_198 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_81_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_81_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_22 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_26 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_81_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_81_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_294 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_296 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_30 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_305 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_81_309 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_320 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_327 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_337 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_81_341 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_81_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_353 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_361 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_369 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_81_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_81_391 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_407 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_41 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_81_410 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_430 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_433 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_437 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_441 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_81_45 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_475 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_482 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_81_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_494 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_81_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_507 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_81_51 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_515 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_81_519 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_523 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_81_532 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_536 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_539 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_547 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_55 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_81_555 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_81_575 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_81_583 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_587 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_590 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_594 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_603 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_607 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_81_611 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_81_627 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_63 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_81_635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_81_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_81_649 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_658 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_81_662 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_81_67 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_81_678 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_682 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_685 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_81_693 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_81_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_81_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_81_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_81_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_81 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_81_84 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_81_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_81_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_81_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_81_929 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_81_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_979 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_981 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_81_984 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_992 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_81_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_10 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_1003 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_82_1007 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_1023 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_1025 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_82_1050 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_1066 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_1068 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_1076 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_82_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_1080 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_1084 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_82_1088 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_1096 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_82_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_82_1134 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_82_1150 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_1158 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_1161 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_1169 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_82_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_82_1205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_1225 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_1233 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_1274 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_1305 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_1309 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_132 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_1324 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_1328 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_1359 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_1363 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_1367 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_14 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_82_140 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_1417 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_1421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_1460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_1464 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_82_1468 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_148 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_82_1500 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_151 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_82_1516 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_1524 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_82_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_82_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_159 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_163 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_167 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_175 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_82_182 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_82_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_82_216 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_24 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_82_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_290 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_82_294 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_82_310 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_82_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_337 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_82_341 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_82_373 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_82_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_82_408 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_420 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_432 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_82_436 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_452 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_465 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_474 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_82_488 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_49 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_504 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_508 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_511 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_515 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_519 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_523 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_53 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_548 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_556 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_569 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_57 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_572 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_584 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_588 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_591 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_608 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_82_61 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_82_614 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_82_646 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_654 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_82_658 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_666 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_685 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_693 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_82_706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_714 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_718 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_82_721 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_82_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_82_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_779 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_786 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_796 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_800 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_82_804 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_81 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_812 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_82_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_83 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_897 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_901 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_82_905 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_921 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_923 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_926 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_930 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_940 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_82_944 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_952 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_956 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_82_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_968 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_972 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_976 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_980 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_83_10 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_83_1032 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_83_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_83_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_83_1083 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_1091 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_1093 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_1096 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_110 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_1100 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_83_1112 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_83_1128 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_83_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_114 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_83_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_1174 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_1178 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_118 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_83_1186 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_83_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_83_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_83_1217 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_83_1224 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_1240 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_1252 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_1260 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_1283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_1300 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_83_1304 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_1310 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_83_1314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_132 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_1333 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_1343 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_1347 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_1367 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_1398 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_14 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_1408 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_1452 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_1456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_1460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_83_1464 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_83_1480 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_1488 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_83_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_151 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_83_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_83_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_162 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_17 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_180 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_83_184 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_83_192 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_196 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_83_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_204 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_83_222 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_83_238 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_248 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_25 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_252 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_83_256 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_83_272 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_83_280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_289 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_297 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_304 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_83_308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_32 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_83_340 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_83_348 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_83_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_41 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_83_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_437 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_83_441 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_83_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_480 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_83_484 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_488 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_49 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_495 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_501 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_507 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_519 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_532 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_540 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_544 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_556 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_56 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_83_564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_83_573 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_58 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_83_581 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_585 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_587 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_590 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_594 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_83_610 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_83_620 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_636 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_644 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_654 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_660 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_662 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_665 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_83_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_680 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_686 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_83_690 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_83_706 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_719 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_726 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_83_730 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_738 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_746 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_83_756 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_76 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_83_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_83_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_80 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_817 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_820 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_828 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_830 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_833 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_857 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_83_861 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_83_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_883 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_887 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_897 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_83_901 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_83_917 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_92 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_921 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_83_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_959 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_83_96 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_966 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_83_970 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_83_986 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_992 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_83_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_10 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_84_1002 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_84_1018 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_1026 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_103 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_84_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_1047 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_1051 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_1055 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_1072 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_1076 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_84_1080 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_84_1096 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_1106 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_111 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_84_1114 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_84_1146 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_84_1154 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_1175 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_1178 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_84_119 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_1190 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_84_1194 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_84_1210 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_1216 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_84_1220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_123 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_84_1232 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_1240 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_84_1248 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_84_1264 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_1272 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_1275 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_1279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_1287 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_1295 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_1299 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_1303 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_1305 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_1366 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_1374 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_1382 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_1402 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_1412 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_84_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_1432 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_1442 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_84_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_148 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_84_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_84_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_155 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_84_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_84_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_84_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_175 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_84_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_84_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_211 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_84_214 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_84_230 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_84_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_26 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_260 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_264 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_84_268 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_84_284 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_290 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_298 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_30 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_308 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_84_312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_316 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_84_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_84_400 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_410 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_423 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_84_427 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_431 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_434 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_438 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_84_44 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_458 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_84_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_84_471 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_477 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_48 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_485 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_495 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_84_51 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_526 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_530 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_84_542 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_55 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_84_552 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_558 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_84_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_84_578 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_84_586 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_84_59 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_590 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_601 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_84_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_609 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_84_612 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_620 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_624 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_639 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_643 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_84_647 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_651 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_653 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_656 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_84_660 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_84_668 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_67 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_672 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_678 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_681 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_84_689 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_84_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_717 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_84_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_721 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_84_725 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_84_741 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_84_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_755 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_757 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_760 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_764 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_84_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_84_80 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_84_804 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_84_812 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_824 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_828 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_84_832 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_84 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_84_848 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_852 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_84_856 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_84_872 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_84_880 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_884 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_84_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_84_921 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_84_929 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_84_945 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_84_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_84_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_84_976 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_990 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_998 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_1012 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_1016 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_85_1020 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_85_1032 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_85_1048 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_1056 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_1076 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_1080 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_85_1084 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_85_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_1130 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_1132 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_1145 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_1154 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_85_1158 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_85_1190 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_85_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_85_1225 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_1233 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_1240 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_85_1255 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_85_127 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_1271 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_1282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_1289 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_85_1293 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_1309 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_1316 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_1318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_1360 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_1367 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_1374 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_1378 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_1380 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_1387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_1395 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_1399 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_1403 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_1409 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_1413 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_1417 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_1431 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_1438 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_85_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_1445 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_1449 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_1453 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_85_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_1489 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_85_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_152 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_156 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_85_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_159 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_85_163 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_85_195 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_85_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_211 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_85_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_85_231 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_239 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_246 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_248 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_251 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_85_260 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_85_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_85_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_85_30 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_322 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_326 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_336 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_85_340 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_348 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_85_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_365 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_368 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_85_376 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_38 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_394 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_85_402 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_418 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_42 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_85_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_85_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_85_476 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_484 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_85_487 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_495 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_503 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_505 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_510 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_541 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_543 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_549 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_555 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_56 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_573 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_579 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_85_583 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_60 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_85_615 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_623 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_627 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_635 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_64 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_647 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_85_671 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_68 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_703 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_707 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_85_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_85_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_748 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_750 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_85_753 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_85_769 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_777 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_85_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_81 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_85_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_823 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_827 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_85_831 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_85 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_863 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_867 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_869 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_872 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_879 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_85_883 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_91 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_915 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_919 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_948 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_85_95 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_85_952 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_85_984 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_992 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_85_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_86_1003 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_1007 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_1015 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_1019 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_1021 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_1040 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_86_1048 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_86_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_1068 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_1071 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_1089 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_1093 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_1097 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_86_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_111 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_86_1110 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_1114 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_1117 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_1121 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_1133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_86_1146 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_86_1162 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_86_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_1189 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_86_1200 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_122 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_86_1232 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_1240 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_1247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_86_1255 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_126 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_1271 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_1274 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_1278 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_1282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_86_1296 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_86_130 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_86_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_1319 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_1322 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_86_1330 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_1334 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_1364 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_1368 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_1372 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_1376 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_86_138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_86_1380 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_1393 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_1397 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_86_1401 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_1407 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_1411 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_86_1423 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_1427 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_1434 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_1438 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_1446 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_86_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_86_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_146 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_86_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_86_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_86_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_86_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_160 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_86_164 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_86_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_86_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_86_187 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_191 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_193 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_86_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_200 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_86_204 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_86_236 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_86_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_86_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_26 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_28 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_86_31 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_86_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_86_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_86_337 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_345 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_361 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_86_365 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_86_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_86_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_395 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_402 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_86_406 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_86_438 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_45 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_86_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_458 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_86_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_467 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_86_470 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_48 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_86_502 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_86_512 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_516 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_86_519 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_585 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_86_589 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_86_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_601 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_612 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_86_616 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_86_648 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_86_664 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_668 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_670 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_688 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_86_692 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_708 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_711 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_715 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_86_719 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_86_735 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_743 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_75 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_751 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_755 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_794 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_86_798 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_814 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_86_827 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_84 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_868 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_86_872 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_86_880 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_86_896 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_86_904 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_908 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_910 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_913 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_917 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_86_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_93 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_86_963 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_97 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_86_995 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_87_10 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_1007 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_1011 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_87_1015 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_1019 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_87_1022 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_87_1030 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_87_1036 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_87_1046 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_87_1054 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_87_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_87_1091 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_87_1123 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_87_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_1140 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_1143 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_87_1151 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_87_116 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_87_1183 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_1191 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_1195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_120 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_87_1203 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_87_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_1217 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_122 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_1225 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_87_1233 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_87_1245 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_87_1284 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_129 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_1300 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_1304 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_1311 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_87_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_1319 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_1323 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_1327 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_87_133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_1331 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_1341 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_1343 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_1346 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_1354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_1358 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_1362 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_1366 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_1368 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_1375 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_1387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_1391 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_87_1395 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_1399 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_14 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_1402 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_1406 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_1410 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_1414 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_1418 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_1425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_1429 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_87_1433 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_1437 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_87_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_1440 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_87_1444 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_87_1476 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_148 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_87_1484 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_1488 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_87_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_150 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_153 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_87_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_87_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_157 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_16 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_161 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_178 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_87_182 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_186 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_19 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_190 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_198 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_87_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_87_218 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_87_234 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_87_242 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_246 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_248 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_87_251 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_87_267 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_87_275 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_87_29 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_295 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_87_299 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_87_331 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_87_347 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_87_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_375 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_382 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_87_386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_87_404 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_87_412 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_87_418 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_87_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_44 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_444 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_448 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_452 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_468 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_478 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_48 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_482 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_87_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_87_517 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_87_52 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_523 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_529 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_87_580 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_586 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_87_590 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_87_606 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_610 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_616 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_87_620 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_636 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_87_645 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_87_653 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_657 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_660 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_664 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_68 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_685 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_689 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_693 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_714 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_726 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_87_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_87_730 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_87_762 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_778 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_87_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_87_81 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_87_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_87_823 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_87_829 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_87_845 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_849 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_85 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_87_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_87_870 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_876 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_88 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_880 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_87_92 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_928 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_932 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_87_936 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_87_944 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_948 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_951 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_87_955 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_968 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_87_972 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_988 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_990 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_1034 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_88_1041 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_1045 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_88_1054 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_88_1062 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_1066 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_88_1069 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_88_1085 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_88_1093 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_1097 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_110 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_88_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_88_1118 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_1132 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_88_1136 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_1152 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_88_1155 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_88_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_118 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_88_1189 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_1199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_88_1203 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_88_122 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_88_1235 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_1250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_1257 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_126 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_88_1261 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_129 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_88_1293 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_1309 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_1317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_1331 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_1335 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_1339 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_88_1343 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_1349 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_1359 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_1363 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_1367 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_1371 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_88_1375 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_88_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_1390 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_1392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_88_1395 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_1403 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_1405 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_88_1408 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_88_1414 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_1418 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_1425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_88_1429 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_143 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_88_1445 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_1453 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_88_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_88_150 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_88_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_88_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_88_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_88_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_161 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_169 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_88_173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_88_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_183 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_88_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_200 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_88_220 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_88_228 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_232 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_235 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_263 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_267 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_88_271 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_28 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_88_303 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_88_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_32 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_334 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_338 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_88_342 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_88_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_88_374 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_88_382 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_386 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_88_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_402 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_414 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_88_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_88_45 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_88_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_88_477 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_88_509 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_88_525 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_529 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_88_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_55 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_88_550 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_556 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_566 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_573 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_577 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_579 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_582 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_88_586 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_88_59 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_590 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_608 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_612 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_643 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_88_651 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_659 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_88_663 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_88_67 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_88_683 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_88_689 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_88_697 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_701 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_71 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_88_717 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_88_733 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_74 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_88_741 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_88_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_88_779 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_88_787 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_88_793 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_88_809 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_813 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_88_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_88_82 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_88_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_896 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_88_900 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_88_916 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_88_924 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_928 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_932 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_936 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_88_944 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_88_952 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_956 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_88_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_88_976 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_88_98 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_980 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_982 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_985 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_88_997 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_89_10 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_100 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_1012 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_1014 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_1021 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_1033 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_1037 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_89_1041 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_89_1057 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_89_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_89_1075 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_1079 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_89_1091 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_89_1107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_1115 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_1117 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_89_1120 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_1140 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_1143 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_1153 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_89_1161 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_89_1177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_118 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_1185 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_1189 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_89_1197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_89_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_89_126 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_89_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_1284 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_89_1288 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_89_1320 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_89_1336 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_1340 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_89_1343 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_1347 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_89_1354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_1364 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_1368 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_89_1372 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_14 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_89_1404 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_89_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_89_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_148 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_89_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_89_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_89_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_89_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_16 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_162 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_168 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_89_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_187 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_190 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_197 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_89_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_211 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_89_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_89_249 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_295 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_299 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_89_303 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_89_335 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_35 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_351 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_89_364 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_372 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_89_375 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_89_39 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_89_407 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_411 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_413 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_89_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_424 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_89_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_444 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_448 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_452 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_491 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_495 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_89_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_89_515 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_523 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_525 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_535 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_89_539 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_89_55 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_89_555 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_572 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_89_575 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_89_591 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_89_606 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_610 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_613 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_623 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_89_627 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_63 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_89_635 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_647 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_89_651 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_89_661 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_665 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_671 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_89_675 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_679 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_682 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_689 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_89_693 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_89_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_718 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_89_726 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_89_758 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_89_774 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_778 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_790 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_792 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_798 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_89_802 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_89_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_89_826 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_830 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_89_833 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_84 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_849 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_89_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_89_88 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_89_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_929 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_933 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_943 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_89_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_89_96 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_89_979 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_89_987 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_991 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_89_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_8_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_8_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_8_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_8_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_8_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_8_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_8_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_8_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_8_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_8_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_8_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_8_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_8_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_8_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_8_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_8_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_8_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_8_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_8_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_8_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_8_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_8_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_8_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_8_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_1027 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_90_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_1037 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_90_1045 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_90_1061 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_1065 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_90_1068 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_90_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_1105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_1109 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_1118 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_1129 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_1133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_1137 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_90_1141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_90_1149 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_90_1155 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_116 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_90_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_90_1189 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_90_1199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_90_1231 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_90_1255 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_90_126 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_90_1271 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_1275 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_1284 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_1291 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_90_1295 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_1311 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_90_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_90_1323 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_1327 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_90_1330 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_90_1346 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_1356 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_90_1360 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_90_1376 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_90_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_90_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_90_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_90_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_90_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_90_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_90_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_90_158 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_90_164 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_90_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_90_182 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_90_190 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_194 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_196 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_90_199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_90_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_90_231 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_90_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_28 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_90_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_32 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_90_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_90_353 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_361 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_90_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_90_373 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_379 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_90_383 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_90_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_90_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_90_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_90_495 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_90_503 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_507 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_514 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_518 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_520 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_90_53 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_536 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_90_539 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_90_547 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_551 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_553 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_556 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_560 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_57 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_60 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_90_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_90_621 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_90_627 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_64 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_90_643 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_90_649 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_90_665 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_90_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_90_708 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_716 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_718 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_90_721 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_90_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_74 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_741 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_749 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_90_756 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_788 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_90_792 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_90_808 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_90_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_82 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_822 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_825 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_90_829 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_90_841 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_86 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_90_873 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_881 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_883 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_90_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_90_90 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_90_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_90_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_992 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_90_995 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_91_10 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_1007 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_91_1011 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_91_1027 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_91_1034 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_91_1050 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_91_1058 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_91_1076 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_91_1108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_1116 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_91_1120 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_91_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_115 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_91_1154 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_1158 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_1165 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_91_1169 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_1187 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_91_1212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_125 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_1276 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_1282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_1285 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_91_129 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_91_1295 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_91_1311 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_1321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_1328 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_133 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_91_1337 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_91_1345 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_91_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_14 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_91_1429 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_146 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_91_1461 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_91_1477 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_91_1485 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_1489 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_91_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_91_153 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_91_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_91_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_169 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_91_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_91_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_204 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_91_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_222 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_91_226 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_230 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_232 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_91_235 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_91_267 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_91_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_33 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_91_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_91_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_91_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_91_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_91_405 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_413 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_420 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_424 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_435 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_91_439 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_91_45 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_91_455 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_459 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_461 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_91_464 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_49 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_91_537 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_543 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_91_547 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_566 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_573 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_625 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_91_63 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_91_633 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_637 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_91_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_91_649 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_91_655 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_659 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_91_663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_67 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_671 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_91_675 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_719 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_726 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_91_730 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_91_762 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_91_770 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_91_790 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_82 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_91_822 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_91_838 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_91_846 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_850 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_860 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_864 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_91_868 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_876 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_884 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_91_894 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_90 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_91_910 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_91_932 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_91_94 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_91_948 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_956 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_958 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_91_961 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_91_977 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_985 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_987 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_92_1001 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_1009 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_92_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_1011 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_1014 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_1018 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_92_1025 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_1033 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_92_1042 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_92_1058 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_92_1068 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_92_1076 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_1080 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_1082 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_92_1085 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_92_1093 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_1097 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_92_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_1110 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_1113 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_1117 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_92_1159 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_1167 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_1182 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_92_1186 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_92_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_92_1210 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_1214 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_92_1217 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_92_1225 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_1231 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_92_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_92_1276 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_1284 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_92_1287 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_92_1303 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_1311 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_92_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_132 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_1331 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_92_1339 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_134 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_92_1371 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_1403 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_1409 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_92_1413 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_92_1429 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_1433 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_1435 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_1442 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_92_1446 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_145 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_92_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_92_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_92_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_92_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_92_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_92_182 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_92_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_214 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_92_218 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_22 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_222 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_225 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_233 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_253 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_92_257 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_267 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_270 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_92_278 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_92_294 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_298 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_302 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_306 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_316 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_32 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_324 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_333 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_92_337 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_92_369 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_373 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_375 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_388 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_92_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_92_40 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_92_424 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_92_440 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_448 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_453 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_469 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_92_473 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_92_505 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_92_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_529 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_56 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_568 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_579 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_585 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_589 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_59 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_593 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_595 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_612 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_92_616 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_620 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_622 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_92_625 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_92_633 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_637 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_639 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_642 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_646 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_653 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_661 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_668 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_670 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_690 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_92_694 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_92_710 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_714 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_716 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_719 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_723 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_734 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_92_738 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_749 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_92_758 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_78 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_92_790 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_92_806 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_814 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_92_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_88 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_92_900 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_92 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_92_932 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_948 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_950 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_96 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_972 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_92_976 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_98 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_984 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_92_991 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_997 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_93_1077 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_1083 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_1093 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_93_1097 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_1113 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_1117 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_93_1121 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_93_1129 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_1133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_93_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_93_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_93_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_93_1215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_93_1229 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_93_1261 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_93_1269 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_1289 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_93_1293 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_93_1309 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_1313 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_1317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_132 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_1321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_93_1330 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_1346 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_93_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_1359 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_93_1367 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_93_1399 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_93_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_1429 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_93_1433 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_93_1465 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_147 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_93_1481 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_1489 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_149 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_93_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_93_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_93_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_93_173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_93_186 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_93_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_93_202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_210 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_93_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_93_231 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_235 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_238 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_248 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_252 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_93_256 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_93_272 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_93_280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_288 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_93_291 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_93_323 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_331 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_333 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_93_336 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_93_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_93_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_373 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_379 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_93_383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_93_415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_423 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_93_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_93_462 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_494 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_93_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_93_50 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_93_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_93_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_578 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_93_58 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_93_583 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_599 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_601 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_93_604 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_93_612 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_616 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_62 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_620 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_93_628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_636 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_64 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_93_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_93_657 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_93_663 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_93_67 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_93_679 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_687 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_691 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_93_699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_707 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_93_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_789 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_93_793 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_93_809 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_813 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_826 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_828 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_831 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_838 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_93_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_850 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_93_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_93_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_93_928 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_936 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_93_939 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_97 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_93_971 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_93_987 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_991 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_93_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_10 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_103 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_94_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_94_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_94_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_94_111 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_94_1134 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_115 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_94_1150 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_94_1160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_1168 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_117 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_94_1176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_94_120 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_94_1208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_1216 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_94_1219 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_94_1227 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_1231 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_94_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_1266 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_94_1270 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_94_128 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_94_1302 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_1310 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_1318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_132 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_1325 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_94_1329 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_94_1337 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_1343 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_94_1371 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_94_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_94_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_1394 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_1398 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_94_140 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_94_1406 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_94_1438 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_94_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_94_150 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_94_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_94_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_94_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_94_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_158 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_161 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_17 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_175 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_94_192 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_94_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_94_224 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_94_240 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_25 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_94_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_94_266 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_274 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_94_289 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_29 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_295 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_94_299 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_94_315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_325 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_33 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_331 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_333 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_336 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_94_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_94_378 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_94_386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_94_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_94_40 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_94_400 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_404 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_406 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_413 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_94_417 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_94_433 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_94_441 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_445 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_94_466 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_48 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_94_482 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_50 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_500 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_504 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_94_508 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_512 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_515 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_519 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_94_53 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_537 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_94_541 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_57 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_94_573 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_94_583 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_59 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_593 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_94_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_601 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_94_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_62 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_94_637 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_653 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_655 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_94_658 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_94_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_74 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_94_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_94_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_94_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_94_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_85 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_850 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_852 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_94_855 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_871 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_875 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_94_883 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_94_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_89 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_94_905 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_913 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_916 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_94_920 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_94_93 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_94_931 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_94_937 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_94_963 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_99 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_94_997 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_1004 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_95_1008 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_1012 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_1016 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_1020 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_103 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_1035 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_1043 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_95_1051 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_95_1059 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_106 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_1063 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_95_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_95_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_1103 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_1113 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_95_1117 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_1133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_95_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_1156 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_1160 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_95_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_1177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_118 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_95_1184 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_95_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_1198 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_1205 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_95_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_95_1243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_1275 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_128 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_95_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_1314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_1317 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_95_132 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_1321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_95_1333 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_95_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_95_1385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_140 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_1417 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_95_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_146 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_95_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_149 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_95_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_95_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_95_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_157 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_168 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_95_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_180 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_184 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_95_188 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_95_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_95_204 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_22 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_222 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_95_226 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_95_258 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_95_274 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_95_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_95_302 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_306 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_309 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_313 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_95_323 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_337 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_95_341 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_95_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_353 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_95_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_95_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_95_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_95_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_476 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_483 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_95_487 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_495 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_95_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_51 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_513 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_95_517 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_95_549 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_95_55 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_95_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_95_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_578 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_581 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_585 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_587 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_59 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_594 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_95_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_614 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_618 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_62 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_95_622 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_643 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_646 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_656 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_665 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_95_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_95_701 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_718 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_95_722 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_730 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_733 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_757 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_76 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_761 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_95_765 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_78 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_95_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_787 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_791 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_795 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_95_803 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_95_835 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_95_843 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_887 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_891 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_95_895 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_901 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_95_909 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_91 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_95_917 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_921 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_95_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_95_933 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_937 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_95_941 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_95_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_961 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_95_965 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_95_981 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_95_99 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_96_1004 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_96_1020 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_96_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_96_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_1043 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_1045 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_1048 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_96_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_96_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_1068 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_1072 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_96_1076 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_96_1086 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_96_1094 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_1098 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_96_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_111 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_96_1134 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_115 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_96_1150 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_1158 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_96_1162 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_1175 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_96_1178 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_96_1210 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_1226 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_1229 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_96_1251 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_96_127 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_1285 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_1289 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_1305 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_96_1309 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_96_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_96_1331 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_1337 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_1341 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_96_1349 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_96_1365 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_1373 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_1377 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_1381 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_96_1405 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_96_1437 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_145 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_1453 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_96_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_149 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_96_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_96_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_96_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_96_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_96_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_182 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_96_186 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_194 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_198 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_96_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_202 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_96_216 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_226 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_96_230 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_238 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_240 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_259 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_96_263 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_96_295 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_32 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_330 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_337 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_96_341 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_96_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_353 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_355 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_96_358 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_374 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_376 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_96_395 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_96_40 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_96_403 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_407 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_409 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_412 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_441 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_445 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_96_449 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_473 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_96_477 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_96_493 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_50 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_96_501 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_511 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_96_515 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_52 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_96_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_55 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_59 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_96_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_96_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_63 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_96_637 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_653 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_655 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_96_658 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_96_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_96_692 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_700 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_723 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_96_727 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_743 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_96_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_779 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_786 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_790 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_96_794 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_96_810 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_814 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_96_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_96_850 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_96_858 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_96_864 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_96_880 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_884 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_96_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_96_963 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_97_10 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_97_1003 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_97_1035 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_1041 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_97_1048 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_1070 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_1084 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_97_109 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_97_1092 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_97_1108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_1116 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_1119 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_1123 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_1134 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_97_1141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_97_1149 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_115 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_1153 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_1160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_1164 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_97_1168 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_1205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_1212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_97_1216 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_97_1232 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_1240 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_1242 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_97_1245 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_1249 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_1251 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_1254 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_1267 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_97_1271 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_97_1287 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_97_129 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_97_1319 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_1323 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_1325 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_1328 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_1332 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_97_1354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_97_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_97_1370 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_97_1378 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_1382 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_1384 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_97_1387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_14 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_97_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_97_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_97_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_151 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_97_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_97_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_158 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_16 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_160 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_97_166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_182 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_97_186 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_19 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_97_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_97_202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_222 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_226 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_23 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_230 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_234 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_254 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_264 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_97_268 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_97_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_290 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_293 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_303 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_97_307 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_97_323 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_327 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_330 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_338 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_97_342 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_368 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_372 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_97_376 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_386 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_393 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_397 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_97_401 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_97_417 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_97_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_97_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_97_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_535 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_539 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_546 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_550 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_97_554 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_97_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_566 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_97_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_60 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_97_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_97_610 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_614 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_97_618 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_97_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_97_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_645 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_652 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_97_656 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_97_67 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_674 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_97_682 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_97_698 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_97_706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_97_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_97_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_97_752 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_756 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_763 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_97_767 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_775 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_777 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_790 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_792 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_809 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_813 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_97_817 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_85 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_97_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_864 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_871 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_97_875 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_89 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_97_891 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_97_899 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_903 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_907 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_97_915 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_97_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_97_93 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_97_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_97_967 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_983 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_97_987 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_10 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_100 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_1003 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_98_1007 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_1015 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_1018 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_1026 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_98_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_1047 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_98_1050 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_1058 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_1062 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_1065 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_98_1073 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_1081 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_1083 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_98_1086 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_1094 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_1096 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_98_1109 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_112 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_98_1141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_115 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_1151 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_1159 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_117 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_1176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_1180 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_1182 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_1185 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_1189 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_1200 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_1210 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_1214 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_98_1218 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_98_1234 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_124 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_98_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_1252 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_1256 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_1274 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_98_1278 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_1286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_1290 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_1294 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_1302 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_1306 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_1310 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_98_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_1323 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_1325 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_1328 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_98_1336 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_98_1368 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_98_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_145 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_98_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_149 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_98_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_153 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_98_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_157 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_16 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_161 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_169 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_187 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_191 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_195 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_98_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_20 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_203 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_210 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_214 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_218 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_222 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_232 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_234 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_246 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_256 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_98_260 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_27 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_98_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_284 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_290 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_294 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_98_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_98_325 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_343 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_98_355 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_371 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_375 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_377 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_380 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_388 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_399 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_403 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_98_411 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_443 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_447 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_466 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_98_470 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_48 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_98_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_494 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_498 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_50 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_506 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_98_510 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_518 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_520 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_523 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_53 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_544 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_98_548 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_568 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_57 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_571 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_588 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_592 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_596 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_61 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_616 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_620 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_624 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_98_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_670 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_683 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_98_687 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_71 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_98_719 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_98_735 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_743 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_98_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_98_779 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_787 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_98_793 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_809 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_813 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_98_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_82 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_828 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_835 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_98_839 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_871 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_885 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_98_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_907 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_98_917 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_98_92 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_935 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_939 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_955 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_98_963 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_971 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_975 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_979 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_983 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_99_1003 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_99_1019 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_99_1027 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_1034 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_99_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_1051 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_99_1055 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_1063 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_99_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_99_1083 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_1091 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_99_1103 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_99_1119 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_99_1127 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_99_1145 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_115 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_99_1153 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_1159 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_99_1163 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_99_1171 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_1175 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_1177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_99_1180 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_1188 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_99_1196 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_1212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_99_1216 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_99_123 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_99_1248 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_99_1264 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_127 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_99_1272 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_1276 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_99_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_1288 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_1291 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_1295 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_1297 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_130 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_1302 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_99_1306 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_99_1322 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_99_1330 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_99_1336 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_99_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_99_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_99_1367 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_1377 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_99_138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_1381 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_99_1395 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_99_1411 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_99_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_1430 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_1433 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_99_1441 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_99_1473 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_1489 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_99_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_99_150 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_99_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_99_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_159 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_99_167 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_183 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_187 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_99_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_223 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_99_233 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_260 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_99_264 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_99_280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_99_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_296 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_300 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_307 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_99_323 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_333 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_99_337 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_99_345 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_351 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_368 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_99_372 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_99_404 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_99_420 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_424 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_434 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_438 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_99_442 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_99_474 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_99_490 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_494 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_99_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_99_535 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_99_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_99_62 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_99_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_99_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_99_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_689 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_691 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_694 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_698 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_708 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_99_715 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_731 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_735 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_745 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_99_749 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_76 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_78 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_99_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_99_799 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_99_819 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_99_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_99_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_99_89 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_99_902 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_906 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_916 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_920 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_99_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_95 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_99_99 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_9_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_9_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_9_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_9_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_9_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_9_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_9_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_9_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_9_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_9_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_9_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_9_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_9_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_9_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_9_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_9_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_9_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_9_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_9_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_9_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_9_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_9_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_9_996 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_0 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_10 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_100 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_101 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_102 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_103 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_104 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_105 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_106 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_107 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_108 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_109 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_11 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_110 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_111 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_112 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_113 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_114 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_115 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_116 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_117 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_118 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_119 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_12 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_120 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_121 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_122 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_123 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_124 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_125 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_126 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_127 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_128 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_129 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_13 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_130 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_131 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_132 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_133 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_134 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_135 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_136 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_137 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_138 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_139 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_14 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_140 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_141 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_142 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_143 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_144 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_145 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_146 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_147 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_148 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_149 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_15 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_150 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_151 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_152 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_153 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_154 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_155 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_156 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_157 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_158 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_159 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_16 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_160 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_161 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_162 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_163 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_164 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_165 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_166 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_167 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_168 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_169 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_17 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_170 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_171 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_172 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_173 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_174 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_175 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_176 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_177 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_178 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_179 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_18 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_180 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_181 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_182 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_183 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_184 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_185 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_186 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_187 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_188 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_189 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_19 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_190 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_191 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_192 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_193 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_194 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_195 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_196 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_197 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_198 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_199 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_2 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_20 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_200 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_201 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_202 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_203 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_204 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_205 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_206 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_207 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_208 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_209 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_21 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_210 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_211 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_212 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_213 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_214 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_215 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_216 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_217 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_218 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_219 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_22 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_220 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_221 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_222 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_223 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_224 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_225 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_226 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_227 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_228 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_229 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_23 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_230 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_231 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_232 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_233 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_234 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_235 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_236 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_237 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_238 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_239 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_24 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_240 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_241 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_242 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_243 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_244 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_245 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_246 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_247 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_248 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_249 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_25 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_250 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_251 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_252 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_253 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_254 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_255 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_256 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_257 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_258 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_259 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_26 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_260 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_261 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_262 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_263 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_264 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_265 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_266 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_267 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_268 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_269 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_27 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_270 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_271 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_272 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_273 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_274 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_275 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_276 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_277 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_278 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_279 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_28 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_280 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_281 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_282 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_283 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_284 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_285 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_286 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_287 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_288 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_289 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_29 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_3 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_30 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_31 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_32 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_33 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_34 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_35 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_36 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_37 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_38 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_39 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_4 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_40 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_41 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_42 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_43 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_44 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_45 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_46 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_47 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_48 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_49 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_5 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_50 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_51 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_52 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_53 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_54 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_55 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_56 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_57 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_58 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_59 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_6 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_60 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_61 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_62 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_63 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_64 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_65 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_66 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_67 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_68 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_69 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_7 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_70 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_71 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_72 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_73 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_74 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_75 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_76 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_77 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_78 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_79 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_8 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_80 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_81 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_82 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_83 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_84 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_85 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_86 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_87 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_88 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_89 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_9 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_90 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_91 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_92 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_93 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_94 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_95 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_96 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_97 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_98 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_99 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1000 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1001 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1002 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1003 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1004 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1005 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1006 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1007 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1008 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1009 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1010 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1011 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1012 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1013 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1014 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1015 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1016 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1018 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1019 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1020 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1021 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1022 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1023 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1025 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1026 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1027 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1029 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1030 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1032 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1033 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1034 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1035 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1036 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1037 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1038 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1040 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1041 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1042 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1043 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1045 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1046 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1047 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1048 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1049 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1050 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1051 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1053 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1054 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1055 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1056 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1057 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1058 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1059 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1061 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1062 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1063 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1065 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1066 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1068 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1069 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1070 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1071 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1072 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1073 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1074 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1075 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1076 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1077 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1078 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1079 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1080 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1081 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1082 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1083 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1084 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1085 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1086 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1088 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1089 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1090 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1091 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1092 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1093 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1094 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1096 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1097 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1098 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1100 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1101 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1103 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1104 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1105 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1106 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1107 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1108 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1109 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1110 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1111 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1112 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1113 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1114 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1115 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1116 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1117 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1118 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1119 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1120 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1121 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1123 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1124 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1125 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1126 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1127 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1128 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1129 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1130 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1132 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1133 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1134 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1136 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1137 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1139 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1140 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1141 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1142 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1143 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1144 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1145 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1146 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1147 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1148 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1149 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1150 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1151 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1152 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1153 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1154 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1155 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1156 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1158 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1159 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1160 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1161 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1162 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1163 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1164 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1165 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1167 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1168 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1169 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1171 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1172 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1174 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1175 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1176 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1177 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1178 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1179 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1180 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1181 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1182 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1183 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1184 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1185 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1186 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1187 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1188 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1189 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1190 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1191 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1193 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1194 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1195 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1196 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1197 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1198 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1199 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1200 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1201 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1203 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1204 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1205 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1207 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1208 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1210 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1211 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1212 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1213 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1214 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1215 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1216 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1217 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1218 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1219 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1220 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1222 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1224 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1225 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1226 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1227 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1228 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1229 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1230 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1231 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1232 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1233 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1234 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1235 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1236 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1238 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1239 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1240 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1242 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1243 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1245 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1246 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1247 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1248 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1249 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1250 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1251 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1252 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1253 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1254 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1255 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1256 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1257 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1258 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1259 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1260 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1261 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1262 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1263 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1264 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1265 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1266 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1267 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1268 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1269 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1270 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1271 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1272 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1274 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1275 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1276 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1278 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1279 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1281 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1282 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1283 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1284 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1285 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1286 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1287 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1288 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1289 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1290 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1291 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1292 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1293 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1294 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1295 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1296 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1297 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1298 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1299 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1300 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1301 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1302 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1303 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1304 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1305 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1306 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1307 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1309 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1310 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1311 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1313 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1314 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1316 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1317 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1318 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1319 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1320 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1321 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1322 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1323 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1324 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1325 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1326 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1327 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1328 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1329 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1330 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1331 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1332 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1333 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1334 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1335 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1336 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1337 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1338 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1339 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1340 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1341 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1342 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1343 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1345 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1346 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1347 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1349 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1350 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1352 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1353 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1354 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1355 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1356 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1357 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1358 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1359 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1360 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1361 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1362 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1363 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1364 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1365 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1366 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1367 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1368 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1369 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1370 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1371 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1372 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1373 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1374 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1375 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1376 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1377 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1378 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1380 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1381 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1382 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1384 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1385 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1387 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1388 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1389 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1390 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1391 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1392 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1393 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1394 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1395 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1396 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1397 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1398 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1399 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1400 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1401 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1402 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1403 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1404 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1405 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1406 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1407 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1408 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1409 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1410 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1411 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1412 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1413 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1414 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1416 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1417 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1418 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1420 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1421 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1423 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1424 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1425 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1426 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1427 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1428 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1429 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1430 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1431 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1432 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1433 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1434 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1435 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1436 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1437 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1438 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1439 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1440 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1441 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1442 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1443 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1444 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1445 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1446 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1447 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1448 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1449 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1451 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1452 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1453 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1455 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1456 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1458 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1459 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1460 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1461 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1462 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1463 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1464 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1465 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1466 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1467 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1468 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1469 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1470 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1471 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1472 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1473 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1474 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1475 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1476 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1477 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1478 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1479 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1480 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1481 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1482 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1483 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1484 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1485 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1487 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1488 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1489 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1491 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1492 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1494 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1495 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1496 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1497 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1498 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1499 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1500 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1501 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1502 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1503 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1504 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1505 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1506 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1507 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1508 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1509 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1510 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1511 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1512 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1513 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1514 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1515 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1516 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1517 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1518 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1519 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1520 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1522 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1523 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1524 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1526 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1527 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1529 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1530 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1531 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1532 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1533 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1534 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1535 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1536 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1537 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1538 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1539 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1540 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1541 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1542 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1543 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1544 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1545 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1546 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1547 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1548 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1549 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1550 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1551 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1552 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1553 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1554 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1555 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1556 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1558 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1559 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1562 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1563 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1565 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1566 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1567 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1568 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1569 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1570 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1571 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1572 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1573 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1574 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1575 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1577 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1578 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1579 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1581 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1582 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1583 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1584 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1585 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1586 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1587 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1588 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1589 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1590 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1591 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1592 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1593 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1594 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1595 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1596 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1597 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1598 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1600 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1601 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1602 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1603 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1604 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1605 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1606 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1607 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1608 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1609 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1610 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1611 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1612 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1613 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1614 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1615 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1616 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1617 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1618 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1619 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1620 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1621 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1622 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1623 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1624 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1625 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1626 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1627 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1628 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1629 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1630 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1631 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1633 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1634 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1636 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1637 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1638 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1639 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1640 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1641 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1642 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1643 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1644 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1645 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1646 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1647 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1648 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1649 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1650 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1651 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1652 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1653 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1654 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1655 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1656 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1657 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1658 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1659 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1660 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1661 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1662 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1663 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1664 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1665 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1666 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1668 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1669 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1671 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1672 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1673 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1674 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1675 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1676 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1677 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1678 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1679 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1680 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1681 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1682 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1683 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1684 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1685 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1686 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1687 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1688 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1689 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1690 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1691 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1692 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1693 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1694 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1695 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1696 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1697 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1698 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1699 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1700 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1701 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1702 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1704 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1705 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1707 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1708 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1709 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1710 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1711 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1712 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1713 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1714 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1715 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1716 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1717 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1718 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1719 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1720 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1721 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1722 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1723 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1724 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1725 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1726 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1727 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1728 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1729 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1730 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1731 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1732 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1733 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1734 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1735 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1736 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1737 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1739 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1740 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1742 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1743 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1744 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1745 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1746 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1747 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1748 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1749 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1750 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1751 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1752 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1753 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1754 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1755 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1756 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1757 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1758 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1759 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1760 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1761 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1762 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1763 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1764 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1765 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1766 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1767 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1768 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1769 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1770 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1771 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1772 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1773 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1774 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1775 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1776 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1777 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1778 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1779 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1780 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1781 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1782 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1783 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1784 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1785 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1786 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1787 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1788 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1789 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1790 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1791 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1792 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1793 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1794 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1795 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1796 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1797 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1798 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1799 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1800 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1801 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1802 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1803 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1804 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1805 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1806 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1807 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1808 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1809 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1810 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1811 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1812 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1813 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1814 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1815 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1816 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1817 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1818 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1819 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1820 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1821 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1822 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1823 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1824 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1825 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1826 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1827 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1828 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1829 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1830 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1831 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1832 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1833 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1834 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1835 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1836 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1837 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1838 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1839 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1840 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1841 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1842 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1843 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1844 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1845 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1846 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1847 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1848 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1849 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1850 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1851 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1852 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1853 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1854 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1855 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1856 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1857 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1858 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1859 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1860 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1861 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1862 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1863 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1864 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1865 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1866 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1867 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1868 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1869 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1870 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1871 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1872 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1873 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1874 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1875 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1876 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1877 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1878 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1879 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1880 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1881 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1882 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1883 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1884 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1885 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1886 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1887 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1888 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1889 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1890 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1891 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1892 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1893 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1894 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1895 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1896 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1897 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1898 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1899 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1900 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1901 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1902 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1903 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1904 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1905 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1906 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1907 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1908 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1909 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1910 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1911 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1912 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1913 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1914 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1915 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1916 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1917 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1918 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1919 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1920 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1921 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1922 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1923 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1924 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1925 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1926 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1927 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1928 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1929 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1930 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1931 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1932 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1933 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1934 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1935 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1936 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1937 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1938 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1939 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1940 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1941 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1942 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1943 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1944 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1945 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1946 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1947 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1948 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1949 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1950 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1951 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1952 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1953 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1954 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1955 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1956 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1957 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1958 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1959 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1960 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1961 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1962 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1963 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1964 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1965 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1966 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1967 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1968 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1969 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1970 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1971 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1972 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1973 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1974 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1975 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1976 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1977 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1978 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1979 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1980 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1981 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1982 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1983 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1984 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1985 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1986 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1987 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1988 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1989 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1990 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1991 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1992 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1993 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1994 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1995 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1996 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1997 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1998 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1999 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2000 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2001 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2002 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2003 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2004 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2005 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2006 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2007 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2008 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2009 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2010 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2011 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2012 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2013 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2014 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2015 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2016 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2017 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2018 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2019 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2020 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2021 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2022 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2023 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2024 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2025 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2026 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2027 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2028 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2029 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2030 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2031 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2032 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2033 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2034 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2035 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2036 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2037 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2038 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2039 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2040 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2041 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2042 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2043 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2044 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2045 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2046 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2047 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2048 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2049 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2050 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2051 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2052 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2053 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2054 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2055 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2056 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2057 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2058 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2059 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2060 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2061 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2062 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2063 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2064 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2065 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2066 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2067 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2068 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2069 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2070 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2071 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2072 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2073 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2074 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2075 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2076 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2077 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2078 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2079 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2080 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2081 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2082 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2083 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2084 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2085 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2086 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2087 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2088 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2089 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2090 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2091 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2092 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2093 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2094 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2095 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2096 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2097 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2098 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2099 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2100 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2101 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2102 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2103 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2104 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2105 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2106 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2107 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2108 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2109 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2110 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2111 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2112 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2113 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2114 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2115 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2116 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2117 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2118 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2119 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2120 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2121 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2122 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2123 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2124 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2125 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2126 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2127 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2128 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2129 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2130 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2131 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2132 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2133 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2134 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2135 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2136 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2137 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2138 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2139 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2140 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2141 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2142 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2143 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2144 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2145 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2146 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2147 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2148 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2149 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2150 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2151 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2152 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2153 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2154 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2155 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2156 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2157 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2158 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2159 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2160 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2161 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2162 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2163 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2164 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2165 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2166 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2167 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2168 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2169 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2170 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2171 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2172 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2173 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2174 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2175 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2176 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2177 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2178 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2179 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2180 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2181 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2182 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2183 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2184 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2185 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2186 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2187 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2188 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2189 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2190 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2191 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2192 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2193 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2194 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2195 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2196 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2197 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2198 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2199 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2200 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2201 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2202 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2203 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2204 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2205 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2206 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2207 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2208 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2209 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2210 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2211 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2212 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2213 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2214 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2215 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2216 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2217 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2218 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2219 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2220 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2221 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2222 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2223 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2224 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2225 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2226 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2227 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2228 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2229 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2230 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2231 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2232 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2233 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2234 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2235 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2236 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2237 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2238 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2239 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2240 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2241 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2242 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2243 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2244 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2245 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2246 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2247 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2248 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2249 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2250 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2251 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2252 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2253 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2254 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2255 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2256 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2257 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2258 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2259 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2260 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2261 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2262 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2263 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2264 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2265 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2266 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2267 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2268 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2269 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2270 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2271 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2272 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2273 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2274 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2275 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2276 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2277 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2278 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2279 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2280 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2281 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2282 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2283 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2284 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2285 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2286 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2287 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2288 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2289 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2290 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2291 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2292 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2293 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2294 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2295 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2296 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2297 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2298 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2299 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2300 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2301 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2302 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2303 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2304 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2305 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2306 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2307 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2308 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2309 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2310 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2311 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2312 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2313 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2314 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2315 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2316 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2317 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2318 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2319 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2320 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2321 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2322 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2323 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2324 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2325 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2326 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2327 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2328 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2329 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2330 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2331 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2332 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2333 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2334 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2335 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2336 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2337 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2338 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2339 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2340 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2341 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2342 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2343 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2344 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2345 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2346 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2347 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2348 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2349 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2350 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2351 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2352 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2353 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2354 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2355 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2356 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2357 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2358 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2359 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2360 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2361 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2362 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2363 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2364 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2365 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2366 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2367 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2368 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2369 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2370 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2371 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2372 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2373 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2374 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2375 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2376 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2377 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2378 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2379 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2380 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2381 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2382 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2383 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2384 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2385 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2386 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2387 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2388 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2389 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2390 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2391 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2392 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2393 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2394 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2395 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2396 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2397 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2398 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2399 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2400 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2401 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2402 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2403 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2404 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2405 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2406 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2407 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2408 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2409 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2410 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2411 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2412 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2413 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2414 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2415 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2416 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2417 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2418 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2419 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2420 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2421 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2422 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2423 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2424 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2425 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2426 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2427 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2428 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2429 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2430 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2431 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2432 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2433 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2434 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2435 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2436 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2437 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2438 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2439 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2440 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2441 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2442 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2443 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2444 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2445 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2446 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2447 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2448 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2449 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2450 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2451 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2452 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2453 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2454 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2455 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2456 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2457 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2458 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2459 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2460 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2461 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2462 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2463 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2464 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2465 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2466 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2467 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2468 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2469 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2470 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2471 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2472 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2473 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2474 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2475 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2476 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2477 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2478 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2479 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2480 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2481 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2482 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2483 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2484 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2485 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2486 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2487 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2488 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2489 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2490 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2491 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2492 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2493 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2494 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2495 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2496 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2497 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2498 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2499 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2500 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2501 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2502 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2503 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2504 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2505 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2506 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2507 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2508 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2509 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2510 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2511 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2512 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2513 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2514 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2515 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2516 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2517 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2518 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2519 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2520 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2521 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2522 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2523 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2524 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2525 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2526 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2527 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2528 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2529 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2530 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2531 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2532 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2533 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2534 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2535 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2536 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2537 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2538 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2539 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2540 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2541 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2542 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2543 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2544 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2545 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2546 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2547 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2548 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2549 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2550 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2551 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2552 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2553 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2554 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2555 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2556 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2557 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2558 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2559 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2560 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2561 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2562 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2563 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2564 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2565 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2566 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2567 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2568 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2569 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2570 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2571 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2572 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2573 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2574 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2575 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2576 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2577 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2578 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2579 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2580 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2581 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2582 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2583 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2584 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2585 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2586 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2587 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2588 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2589 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2590 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2591 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2592 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2593 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2594 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2595 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2596 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2597 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2598 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2599 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2600 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2601 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2602 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2603 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2604 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2605 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2606 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2607 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2608 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2609 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2610 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2611 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2612 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2613 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2614 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2615 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2616 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2617 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2618 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2619 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2620 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2621 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2622 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2623 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2624 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2625 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2626 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2627 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2628 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2629 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2630 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2631 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2632 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2633 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2634 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2635 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2636 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2637 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2638 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2639 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2640 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2641 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2642 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2643 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2644 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2645 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2646 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2647 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2648 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2649 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2650 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2651 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2652 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2653 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2654 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2655 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2656 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2657 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2658 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2659 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2660 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2661 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2662 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2663 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2664 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2665 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2666 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2667 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2668 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2669 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2670 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2671 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2672 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2673 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2674 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2675 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2676 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2677 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2678 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2679 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2680 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2681 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2682 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2683 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2684 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2685 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2686 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2687 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2688 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2689 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2690 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2691 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2692 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2693 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2694 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2695 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2696 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2697 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2698 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2699 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2700 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2701 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2702 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2703 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2704 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2705 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2706 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2707 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2708 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2709 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2710 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2711 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2712 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2713 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2714 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2715 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2716 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2717 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2718 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2719 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2720 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2721 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2722 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2723 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2724 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2725 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2726 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2727 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2728 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2729 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2730 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2731 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2732 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2733 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2734 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2735 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2736 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2737 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2738 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2739 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2740 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2741 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2742 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2743 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2744 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2745 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2746 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2747 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2748 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2749 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2750 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2751 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2752 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2753 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2754 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2755 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2756 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2757 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2758 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2759 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2760 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2761 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2762 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2763 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2764 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2765 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2766 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2767 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2768 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2769 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2770 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2771 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2772 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2773 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2774 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2775 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2776 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2777 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2778 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2779 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2780 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2781 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2782 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2783 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2784 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2785 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2786 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2787 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2788 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2789 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2790 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2791 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2792 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2793 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2794 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2795 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2796 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2797 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2798 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2799 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2800 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2801 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2802 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2803 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2804 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2805 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2806 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2807 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2808 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2809 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2810 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2811 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2812 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2813 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2814 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2815 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2816 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2817 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2818 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2819 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2820 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2821 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2822 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2823 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2824 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2825 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2826 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2827 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2828 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2829 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2830 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2831 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2832 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2833 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2834 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2835 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2836 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2837 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2838 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2839 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2840 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2841 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2842 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2843 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2844 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2845 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2846 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2847 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2848 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2849 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2850 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2851 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2852 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2853 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2854 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2855 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2856 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2857 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2858 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2859 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2860 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2861 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2862 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2863 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2864 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2865 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2866 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2867 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2868 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2869 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2870 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2871 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2872 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2873 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2874 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2875 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2876 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2877 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2878 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2879 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2880 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2881 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2882 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2883 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2884 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2885 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2886 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2887 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2888 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2889 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2890 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2891 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2892 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2893 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2894 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2895 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2896 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2897 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2898 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2899 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_290 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2900 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2901 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2902 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2903 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2904 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2905 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2906 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2907 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2908 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2909 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_291 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2910 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2911 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2912 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2913 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2914 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2915 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2916 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2917 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2918 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2919 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_292 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2920 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2921 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2922 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2923 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2924 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2925 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2926 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2927 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2928 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2929 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_293 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2930 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2931 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2932 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2933 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2934 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2935 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2936 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2937 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2938 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2939 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_294 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2940 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2941 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2942 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2943 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2944 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2945 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2946 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2947 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2948 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2949 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_295 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2950 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2951 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2952 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2953 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2954 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2955 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2956 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2957 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2958 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2959 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_296 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2960 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2961 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2962 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2963 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2964 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2965 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2966 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2967 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2968 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2969 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_297 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2970 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2971 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2972 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2973 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2974 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2975 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2976 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2977 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2978 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2979 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_298 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2980 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2981 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2982 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2983 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2984 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2985 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2986 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2987 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2988 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2989 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_299 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2990 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2991 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2992 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2993 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2994 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2995 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2996 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2997 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2998 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2999 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_300 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3000 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3001 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3002 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3003 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3004 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3005 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3006 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3007 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3008 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3009 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_301 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3010 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3011 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3012 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3013 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3014 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3015 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3016 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3017 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3018 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3019 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_302 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3020 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3021 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3022 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3023 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3024 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3025 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3026 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3027 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3028 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3029 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_303 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3030 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3031 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3032 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3033 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3034 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3035 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3036 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3037 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3038 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3039 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_304 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3040 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3041 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3042 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3043 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3044 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3045 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3046 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3047 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3048 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3049 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_305 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3050 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3051 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3052 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3053 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3054 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3055 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3056 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3057 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3058 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3059 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_306 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3060 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3061 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3062 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3063 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3064 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3065 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3066 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3067 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3068 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3069 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_307 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3070 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3071 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3072 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3073 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3074 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3075 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3076 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3077 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3078 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3079 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_308 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3080 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3081 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3082 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3083 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3084 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3085 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3086 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3087 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3088 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3089 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_309 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3090 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3091 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3092 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3093 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3094 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3095 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3096 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3097 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3098 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3099 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_310 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3100 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3101 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3102 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3103 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3104 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3105 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3106 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3107 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3108 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3109 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_311 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3110 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3111 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3112 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3113 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3114 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3115 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3116 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3117 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3118 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3119 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_312 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3120 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3121 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3122 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3123 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3124 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3125 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3126 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3127 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3128 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3129 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_313 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3130 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3131 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3132 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3133 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3134 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3135 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3136 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3137 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3138 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3139 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_314 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3140 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3141 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3142 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3143 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3144 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3145 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3146 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3147 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3148 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3149 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_315 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3150 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3151 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3152 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3153 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3154 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3155 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3156 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3157 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3158 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3159 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_316 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3160 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3161 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3162 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3163 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3164 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3165 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3166 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3167 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3168 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3169 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_317 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3170 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3171 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3172 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3173 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3174 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3175 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3176 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3177 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3178 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3179 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_318 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3180 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3181 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3182 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3183 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3184 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3185 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3186 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3187 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3188 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3189 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_319 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3190 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3191 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3192 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3193 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3194 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3195 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3196 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3197 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3198 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3199 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_320 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3200 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3201 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3202 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3203 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3204 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3205 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3206 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3207 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3208 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3209 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_321 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3210 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3211 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3212 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3213 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3214 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3215 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3216 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3217 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3218 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3219 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_322 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3220 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3221 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3222 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3223 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3224 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3225 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3226 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3227 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3228 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3229 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_323 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3230 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3231 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3232 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3233 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3234 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3235 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3236 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3237 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3238 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3239 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_324 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3240 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3241 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3242 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3243 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3244 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3245 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3246 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3247 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3248 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3249 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_325 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3250 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3251 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3252 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3253 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3254 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3255 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3256 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3257 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3258 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3259 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_326 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3260 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3261 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3262 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3263 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3264 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3265 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3266 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3267 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3268 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3269 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_327 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3270 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3271 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3272 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3273 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3274 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3275 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3276 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3277 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3278 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3279 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_328 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3280 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3281 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3282 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3283 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3284 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3285 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3286 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3287 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3288 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3289 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_329 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3290 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3291 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3292 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3293 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3294 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3295 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3296 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3297 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3298 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3299 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_330 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3300 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3301 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3302 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3303 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3304 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3305 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3306 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3307 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3308 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3309 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_331 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3310 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3311 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3312 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3313 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3314 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3315 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3316 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3317 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3318 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3319 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_332 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3320 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3321 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3322 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3323 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3324 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3325 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3326 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3327 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3328 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3329 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_333 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3330 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3331 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3332 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3333 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3334 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3335 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3336 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3337 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3338 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3339 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_334 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3340 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3341 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3342 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3343 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3344 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3345 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3346 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3347 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3348 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3349 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_335 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3350 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3351 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3352 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3353 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3354 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3355 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3356 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3357 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3358 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3359 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_336 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3360 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3361 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3362 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3363 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3364 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3365 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3366 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3367 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3368 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3369 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_337 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3370 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3371 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3372 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3373 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3374 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3375 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3376 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3377 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3378 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3379 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_338 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3380 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3381 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3382 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3383 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3384 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3385 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3386 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3387 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3388 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3389 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_339 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3390 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3391 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3392 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3393 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3394 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3395 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3396 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3397 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3398 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3399 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_340 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3400 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3401 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3402 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3403 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3404 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3405 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3406 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3407 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3408 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3409 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_341 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3410 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3411 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3412 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3413 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3414 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3415 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3416 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3417 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3418 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3419 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_342 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3420 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3421 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3422 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3423 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3424 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3425 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3426 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3427 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3428 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3429 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_343 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3430 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3431 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3432 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3433 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3434 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3435 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3436 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3437 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3438 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3439 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_344 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3440 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3441 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3442 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3443 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3444 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3445 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3446 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3447 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3448 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3449 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_345 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3450 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3451 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3452 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3453 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3454 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3455 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3456 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3457 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3458 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3459 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_346 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3460 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3461 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3462 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3463 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3464 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3465 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3466 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3467 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3468 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3469 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_347 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3470 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3471 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3472 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3473 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3474 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3475 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3476 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3477 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3478 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3479 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_348 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3480 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3481 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3482 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3483 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3484 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3485 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3486 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3487 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3488 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3489 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_349 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3490 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3491 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3492 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3493 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3494 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3495 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3496 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3497 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3498 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3499 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_350 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3500 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3501 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3502 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3503 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3504 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3505 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3506 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3507 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3508 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3509 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_351 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3510 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3511 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3512 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3513 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3514 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3515 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3516 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3517 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3518 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3519 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_352 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3520 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3521 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3522 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3523 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3524 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3525 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_353 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_354 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_355 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_356 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_357 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_358 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_359 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_360 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_361 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_362 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_363 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_364 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_365 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_366 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_367 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_368 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_369 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_370 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_371 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_372 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_373 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_374 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_375 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_376 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_377 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_378 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_379 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_380 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_381 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_382 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_383 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_384 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_385 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_386 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_387 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_388 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_389 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_390 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_391 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_392 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_393 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_394 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_395 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_396 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_397 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_398 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_399 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_400 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_401 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_402 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_403 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_404 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_405 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_406 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_407 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_408 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_409 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_410 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_411 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_412 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_413 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_414 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_415 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_416 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_417 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_418 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_419 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_420 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_421 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_422 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_423 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_424 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_425 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_426 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_427 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_428 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_429 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_430 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_431 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_432 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_433 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_434 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_435 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_436 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_437 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_438 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_439 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_440 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_441 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_442 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_443 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_444 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_445 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_446 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_447 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_448 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_449 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_450 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_451 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_452 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_453 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_454 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_455 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_456 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_457 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_458 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_459 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_460 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_461 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_462 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_463 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_464 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_465 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_466 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_467 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_468 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_469 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_470 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_471 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_472 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_473 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_474 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_475 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_476 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_477 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_478 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_479 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_480 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_481 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_482 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_483 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_484 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_485 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_486 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_487 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_488 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_489 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_490 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_491 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_492 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_493 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_494 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_495 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_496 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_497 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_498 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_499 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_500 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_501 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_502 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_503 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_504 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_505 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_506 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_507 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_508 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_509 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_510 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_511 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_512 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_513 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_514 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_515 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_516 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_517 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_518 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_519 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_520 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_521 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_522 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_523 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_524 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_525 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_526 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_527 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_528 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_529 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_530 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_531 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_532 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_533 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_534 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_535 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_536 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_537 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_538 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_539 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_540 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_541 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_542 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_543 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_544 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_545 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_546 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_547 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_548 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_549 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_550 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_551 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_552 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_553 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_554 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_555 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_556 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_557 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_558 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_559 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_560 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_561 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_562 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_563 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_564 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_565 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_566 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_567 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_568 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_569 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_570 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_571 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_572 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_573 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_574 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_575 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_576 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_577 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_578 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_579 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_580 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_581 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_582 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_583 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_584 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_585 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_586 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_587 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_588 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_589 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_590 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_591 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_592 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_593 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_594 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_595 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_596 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_597 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_598 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_599 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_600 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_601 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_602 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_603 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_604 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_605 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_606 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_607 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_608 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_609 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_610 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_611 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_612 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_613 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_614 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_615 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_616 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_617 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_618 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_619 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_620 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_621 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_622 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_623 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_624 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_625 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_626 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_627 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_628 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_629 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_630 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_631 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_632 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_633 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_634 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_635 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_636 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_637 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_638 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_639 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_640 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_641 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_642 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_643 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_644 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_645 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_646 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_647 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_648 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_649 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_650 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_651 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_652 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_653 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_654 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_655 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_656 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_657 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_658 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_659 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_660 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_661 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_662 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_663 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_664 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_665 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_666 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_667 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_668 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_669 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_670 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_671 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_672 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_673 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_674 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_675 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_676 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_677 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_678 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_679 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_680 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_681 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_682 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_683 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_684 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_685 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_686 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_687 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_688 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_689 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_690 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_691 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_692 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_693 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_694 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_695 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_696 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_697 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_698 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_699 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_700 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_701 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_702 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_703 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_704 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_705 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_706 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_707 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_708 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_709 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_710 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_711 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_712 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_713 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_714 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_715 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_716 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_717 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_718 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_719 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_720 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_721 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_722 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_723 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_724 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_725 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_726 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_727 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_728 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_729 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_730 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_731 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_732 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_733 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_734 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_735 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_736 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_737 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_738 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_739 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_740 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_741 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_742 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_743 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_744 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_745 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_746 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_747 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_748 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_749 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_750 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_751 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_752 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_753 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_754 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_755 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_756 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_757 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_758 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_759 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_760 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_761 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_762 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_763 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_764 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_765 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_766 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_767 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_768 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_769 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_770 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_771 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_772 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_773 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_774 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_775 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_776 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_777 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_778 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_779 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_780 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_781 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_782 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_783 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_784 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_785 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_786 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_787 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_788 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_789 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_790 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_791 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_792 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_793 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_794 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_795 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_796 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_797 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_798 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_799 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_800 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_801 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_802 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_803 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_804 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_805 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_806 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_807 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_808 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_809 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_810 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_811 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_812 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_813 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_814 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_815 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_816 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_817 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_818 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_819 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_820 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_821 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_822 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_823 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_824 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_825 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_826 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_827 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_828 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_829 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_830 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_831 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_832 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_833 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_834 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_835 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_836 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_837 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_838 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_839 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_840 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_841 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_842 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_843 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_844 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_845 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_846 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_847 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_848 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_849 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_850 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_851 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_852 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_853 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_854 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_855 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_856 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_857 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_858 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_859 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_860 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_861 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_862 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_863 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_864 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_865 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_866 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_867 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_868 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_869 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_870 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_871 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_872 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_873 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_874 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_875 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_876 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_877 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_878 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_879 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_880 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_881 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_882 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_883 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_884 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_885 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_886 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_887 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_888 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_889 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_890 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_891 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_892 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_893 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_894 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_895 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_896 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_897 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_898 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_899 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_900 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_901 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_902 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_903 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_904 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_905 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_906 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_907 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_908 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_909 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_910 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_911 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_912 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_913 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_914 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_915 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_916 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_917 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_918 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_919 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_920 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_921 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_922 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_923 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_924 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_925 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_926 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_927 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_928 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_929 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_930 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_931 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_932 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_933 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_934 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_935 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_936 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_937 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_938 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_939 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_940 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_941 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_942 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_943 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_944 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_945 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_946 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_947 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_948 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_949 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_950 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_951 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_952 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_953 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_954 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_955 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_956 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_957 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_958 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_959 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_960 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_961 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_962 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_963 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_964 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_965 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_966 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_967 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_968 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_969 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_970 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_971 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_972 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_973 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_974 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_975 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_976 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_977 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_978 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_979 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_980 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_981 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_982 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_983 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_984 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_985 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_986 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_987 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_988 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_989 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_990 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_991 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_992 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_993 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_994 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_995 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_996 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_997 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_998 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_999 ();
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4553_ (.I(net26),
    .ZN(net13));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4554_ (.I(\as2650.ins_reg[1] ),
    .Z(_4135_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4555_ (.I(_4135_),
    .Z(_4136_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4556_ (.I(_4136_),
    .Z(_4137_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4557_ (.I(\as2650.ins_reg[0] ),
    .Z(_4138_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _4558_ (.I(_4138_),
    .Z(_4139_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _4559_ (.A1(_4139_),
    .A2(_4135_),
    .ZN(_4140_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4560_ (.I(_4140_),
    .Z(_4141_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4561_ (.I(_4141_),
    .Z(_4142_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4562_ (.I(_4142_),
    .Z(_4143_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _4563_ (.I(\as2650.psl[4] ),
    .Z(_4144_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4564_ (.I(_4144_),
    .Z(_4145_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4565_ (.I(_4145_),
    .Z(_4146_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4566_ (.I(_4146_),
    .Z(_4147_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4567_ (.I(_4147_),
    .Z(_4148_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4568_ (.I(_4148_),
    .Z(_4149_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4569_ (.I(_4149_),
    .ZN(_4150_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _4570_ (.A1(\as2650.halted ),
    .A2(net5),
    .ZN(_4151_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4571_ (.I(_4151_),
    .Z(_4152_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4572_ (.A1(_4150_),
    .A2(_4152_),
    .ZN(_4153_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _4573_ (.A1(_4143_),
    .A2(_4153_),
    .ZN(_4154_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4574_ (.I(\as2650.ins_reg[4] ),
    .Z(_4155_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4575_ (.I(_4155_),
    .Z(_4156_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4576_ (.I(_4156_),
    .Z(_4157_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4577_ (.I(\as2650.ins_reg[6] ),
    .Z(_4158_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4578_ (.I(_4158_),
    .Z(_4159_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4579_ (.I(_4159_),
    .Z(_4160_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _4580_ (.A1(_4157_),
    .A2(_4160_),
    .ZN(_4161_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4581_ (.I(\as2650.ins_reg[3] ),
    .Z(_4162_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_4 _4582_ (.A1(\as2650.cycle[7] ),
    .A2(\as2650.cycle[6] ),
    .A3(\as2650.cycle[5] ),
    .A4(\as2650.cycle[4] ),
    .ZN(_4163_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4583_ (.I(\as2650.cycle[2] ),
    .Z(_4164_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4584_ (.A1(\as2650.cycle[3] ),
    .A2(_4164_),
    .ZN(_4165_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4585_ (.I(_4165_),
    .Z(_4166_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _4586_ (.A1(_4163_),
    .A2(_4166_),
    .ZN(_4167_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4587_ (.I(\as2650.cycle[0] ),
    .ZN(_4168_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4588_ (.A1(\as2650.cycle[1] ),
    .A2(_4168_),
    .ZN(_4169_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4589_ (.A1(_4167_),
    .A2(_4169_),
    .ZN(_4170_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4590_ (.A1(_4162_),
    .A2(_4170_),
    .ZN(_4171_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _4591_ (.I(_4163_),
    .Z(_4172_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4592_ (.I(\as2650.cycle[1] ),
    .ZN(_4173_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _4593_ (.I(_4173_),
    .Z(_4174_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _4594_ (.A1(_4174_),
    .A2(_4168_),
    .ZN(_4175_));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _4595_ (.A1(_4172_),
    .A2(_4166_),
    .A3(_4175_),
    .Z(_4176_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4596_ (.I(\as2650.ins_reg[7] ),
    .Z(_4177_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4597_ (.I(_4177_),
    .Z(_4178_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4598_ (.I(_4178_),
    .ZN(_4179_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4599_ (.I(\as2650.ins_reg[2] ),
    .Z(_4180_));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _4600_ (.I(_4180_),
    .ZN(_4181_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4601_ (.I(\as2650.ins_reg[5] ),
    .Z(_4182_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4602_ (.I(_4182_),
    .Z(_4183_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _4603_ (.A1(_4155_),
    .A2(_4183_),
    .Z(_4184_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _4604_ (.A1(_4181_),
    .A2(_4184_),
    .Z(_4185_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4605_ (.A1(_4179_),
    .A2(_4185_),
    .ZN(_4186_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _4606_ (.A1(\as2650.ins_reg[3] ),
    .A2(_4186_),
    .ZN(_4187_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4607_ (.A1(_4176_),
    .A2(_4187_),
    .ZN(_4188_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4608_ (.A1(_4161_),
    .A2(_4171_),
    .B(_4188_),
    .ZN(_4189_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _4609_ (.A1(\as2650.ins_reg[2] ),
    .A2(\as2650.ins_reg[3] ),
    .ZN(_4190_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4610_ (.I(_4190_),
    .Z(_4191_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4611_ (.I(_4183_),
    .Z(_4192_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4612_ (.A1(_4158_),
    .A2(_4177_),
    .ZN(_4193_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_2 _4613_ (.A1(_4156_),
    .A2(_4192_),
    .A3(_4193_),
    .ZN(_4194_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _4614_ (.A1(_4191_),
    .A2(_4194_),
    .Z(_4195_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _4615_ (.I(_4138_),
    .Z(_4196_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4616_ (.I(_4196_),
    .Z(_4197_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _4617_ (.A1(_4197_),
    .A2(_4135_),
    .Z(_4198_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4618_ (.I(_4198_),
    .Z(_4199_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4619_ (.I(\as2650.halted ),
    .Z(_4200_));
 gf180mcu_fd_sc_mcu7t5v0__inv_2 _4620_ (.I(_4200_),
    .ZN(_4201_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4621_ (.I(net5),
    .Z(_4202_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4622_ (.I(_4202_),
    .ZN(_4203_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _4623_ (.A1(_4201_),
    .A2(_4203_),
    .ZN(_4204_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4624_ (.A1(_4149_),
    .A2(_4204_),
    .ZN(_4205_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _4625_ (.A1(_4199_),
    .A2(_4205_),
    .ZN(_4206_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _4626_ (.A1(_4163_),
    .A2(_4165_),
    .Z(_4207_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4627_ (.I(\as2650.cycle[0] ),
    .Z(_4208_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4628_ (.A1(_4173_),
    .A2(_4208_),
    .ZN(_4209_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4629_ (.A1(_4207_),
    .A2(_4209_),
    .ZN(_4210_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _4630_ (.I(_4210_),
    .Z(_4211_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4631_ (.A1(_4206_),
    .A2(_4211_),
    .ZN(_4212_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4632_ (.A1(_4195_),
    .A2(_4212_),
    .ZN(_4213_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4633_ (.I(_4162_),
    .Z(_4214_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4634_ (.I(_4181_),
    .Z(_4215_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _4635_ (.A1(\as2650.ins_reg[4] ),
    .A2(\as2650.ins_reg[6] ),
    .A3(\as2650.ins_reg[7] ),
    .ZN(_4216_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4636_ (.A1(_4182_),
    .A2(_4216_),
    .ZN(_4217_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4637_ (.I(_4217_),
    .Z(_4218_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _4638_ (.A1(_4215_),
    .A2(_4218_),
    .ZN(_4219_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _4639_ (.A1(_4214_),
    .A2(_4219_),
    .ZN(_4220_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4640_ (.A1(_4212_),
    .A2(_4220_),
    .ZN(_4221_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4641_ (.I(_4221_),
    .Z(_4222_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4642_ (.I(_4162_),
    .Z(_4223_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4643_ (.I(_4156_),
    .Z(_4224_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4644_ (.A1(_4159_),
    .A2(_4179_),
    .ZN(_4225_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4645_ (.A1(_4192_),
    .A2(_4225_),
    .ZN(_4226_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _4646_ (.A1(_4181_),
    .A2(_4224_),
    .A3(_4226_),
    .ZN(_4227_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4647_ (.A1(_4223_),
    .A2(_4227_),
    .ZN(_4228_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4648_ (.A1(_4212_),
    .A2(_4228_),
    .ZN(_4229_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4649_ (.I(_4229_),
    .Z(_4230_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4650_ (.I(_4230_),
    .Z(_4231_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4651_ (.I(_4224_),
    .Z(_4232_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _4652_ (.I(_4232_),
    .Z(_4233_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4653_ (.I(\as2650.cycle[7] ),
    .ZN(_4234_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4654_ (.I(_4234_),
    .Z(_4235_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4655_ (.A1(_4173_),
    .A2(\as2650.cycle[0] ),
    .ZN(_4236_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4656_ (.I(_4236_),
    .Z(_4237_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4657_ (.I(\as2650.cycle[6] ),
    .Z(_4238_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4658_ (.A1(\as2650.cycle[5] ),
    .A2(\as2650.cycle[4] ),
    .ZN(_4239_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _4659_ (.A1(_4238_),
    .A2(_4239_),
    .A3(_4165_),
    .ZN(_4240_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _4660_ (.A1(_4237_),
    .A2(_4240_),
    .ZN(_4241_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _4661_ (.A1(_4235_),
    .A2(_4241_),
    .ZN(_4242_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4662_ (.I(\as2650.idx_ctrl[1] ),
    .Z(_4243_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4663_ (.I(\as2650.idx_ctrl[0] ),
    .Z(_4244_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4664_ (.A1(_4243_),
    .A2(_4244_),
    .ZN(_4245_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _4665_ (.I(_4245_),
    .Z(_4246_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_4 _4666_ (.A1(_4233_),
    .A2(_4206_),
    .A3(_4242_),
    .A4(_4246_),
    .ZN(_4247_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4667_ (.I(_4149_),
    .Z(_4248_));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _4668_ (.I(\as2650.ins_reg[4] ),
    .ZN(_4249_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4669_ (.I(_4249_),
    .Z(_4250_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4670_ (.I(\as2650.cycle[3] ),
    .ZN(_4251_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4671_ (.A1(\as2650.cycle[1] ),
    .A2(\as2650.cycle[0] ),
    .ZN(_4252_));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _4672_ (.A1(_4251_),
    .A2(\as2650.cycle[2] ),
    .A3(_4252_),
    .Z(_4253_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4673_ (.A1(_4163_),
    .A2(_4253_),
    .ZN(_4254_));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _4674_ (.I(\as2650.ins_reg[3] ),
    .ZN(_4255_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _4675_ (.A1(_4181_),
    .A2(_4255_),
    .ZN(_4256_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4676_ (.I(_4256_),
    .Z(_4257_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _4677_ (.A1(\as2650.ins_reg[5] ),
    .A2(_4158_),
    .A3(_4177_),
    .ZN(_4258_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _4678_ (.A1(_4198_),
    .A2(_4257_),
    .A3(_4245_),
    .A4(_4258_),
    .ZN(_4259_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _4679_ (.A1(_4254_),
    .A2(_4259_),
    .ZN(_4260_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _4680_ (.A1(_4250_),
    .A2(_4151_),
    .A3(_4260_),
    .ZN(_4261_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4681_ (.A1(_4248_),
    .A2(_4261_),
    .ZN(_4262_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_2 _4682_ (.A1(_4235_),
    .A2(_4236_),
    .A3(_4240_),
    .ZN(_4263_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4683_ (.I(\as2650.addr_buff[6] ),
    .Z(_4264_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4684_ (.I(\as2650.addr_buff[5] ),
    .Z(_4265_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4685_ (.A1(_4264_),
    .A2(_4265_),
    .ZN(_4266_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4686_ (.A1(\as2650.addr_buff[7] ),
    .A2(_4266_),
    .ZN(_4267_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _4687_ (.A1(_4263_),
    .A2(_4267_),
    .ZN(_4268_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_2 _4688_ (.A1(_4233_),
    .A2(_4206_),
    .A3(_4268_),
    .ZN(_4269_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _4689_ (.A1(_4247_),
    .A2(_4262_),
    .A3(_4269_),
    .ZN(_4270_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _4690_ (.A1(_4213_),
    .A2(_4222_),
    .A3(_4231_),
    .A4(_4270_),
    .ZN(_4271_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _4691_ (.A1(_4154_),
    .A2(_4189_),
    .B(_4271_),
    .ZN(_4272_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4692_ (.A1(_4137_),
    .A2(_4272_),
    .ZN(_4273_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4693_ (.I(_4273_),
    .Z(_4274_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4694_ (.I(_4274_),
    .ZN(_4275_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _4695_ (.I(_4262_),
    .Z(_4276_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4696_ (.I(_4192_),
    .Z(_4277_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _4697_ (.A1(_4159_),
    .A2(_4178_),
    .ZN(_4278_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4698_ (.A1(_4277_),
    .A2(_4278_),
    .ZN(_4279_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _4699_ (.A1(_4138_),
    .A2(\as2650.ins_reg[1] ),
    .Z(_4280_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _4700_ (.I0(\as2650.r123[2][0] ),
    .I1(\as2650.r123_2[2][0] ),
    .S(_4147_),
    .Z(_4281_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4701_ (.A1(_4280_),
    .A2(_4281_),
    .ZN(_4282_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4702_ (.I(_4282_),
    .Z(_4283_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4703_ (.I(\as2650.r0[0] ),
    .Z(_4284_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4704_ (.I(_4284_),
    .Z(_4285_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _4705_ (.A1(_4138_),
    .A2(_4135_),
    .Z(_4286_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _4706_ (.I0(\as2650.r123[1][0] ),
    .I1(\as2650.r123[0][0] ),
    .I2(\as2650.r123_2[1][0] ),
    .I3(\as2650.r123_2[0][0] ),
    .S0(\as2650.ins_reg[0] ),
    .S1(_4146_),
    .Z(_4287_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _4707_ (.A1(_4285_),
    .A2(_4140_),
    .B1(_4286_),
    .B2(_4287_),
    .ZN(_4288_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4708_ (.I(_4288_),
    .Z(_4289_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _4709_ (.A1(_4190_),
    .A2(_4283_),
    .A3(_4289_),
    .ZN(_4290_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4710_ (.I(\as2650.holding_reg[0] ),
    .Z(_4291_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4711_ (.A1(_4291_),
    .A2(_4190_),
    .ZN(_4292_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4712_ (.I(_4292_),
    .ZN(_4293_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4713_ (.I(_4285_),
    .Z(_4294_));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _4714_ (.I(_4294_),
    .ZN(_4295_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4715_ (.A1(_4295_),
    .A2(_4198_),
    .ZN(_4296_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4716_ (.I(_4280_),
    .Z(_4297_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4717_ (.I(_4297_),
    .Z(_4298_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _4718_ (.A1(_4298_),
    .A2(_4281_),
    .Z(_4299_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4719_ (.I(_4286_),
    .Z(_4300_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _4720_ (.A1(_4300_),
    .A2(_4287_),
    .Z(_4301_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_2 _4721_ (.A1(_4296_),
    .A2(_4299_),
    .A3(_4301_),
    .B(_4291_),
    .ZN(_4302_));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _4722_ (.A1(_4290_),
    .A2(_4293_),
    .A3(_4302_),
    .Z(_4303_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _4723_ (.A1(_4283_),
    .A2(_4289_),
    .Z(_4304_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4724_ (.I(_4283_),
    .Z(_4305_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4725_ (.I(_4289_),
    .Z(_4306_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4726_ (.I(\as2650.holding_reg[0] ),
    .ZN(_4307_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _4727_ (.A1(_4305_),
    .A2(_4306_),
    .B(_4307_),
    .ZN(_4308_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _4728_ (.A1(_4291_),
    .A2(_4256_),
    .ZN(_4309_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_4 _4729_ (.A1(_4256_),
    .A2(_4304_),
    .B(_4308_),
    .C(_4309_),
    .ZN(_4310_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _4730_ (.A1(_4303_),
    .A2(_4310_),
    .ZN(_4311_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4731_ (.I(_4183_),
    .Z(_4312_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4732_ (.A1(_4159_),
    .A2(_4179_),
    .ZN(_4313_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4733_ (.I(_4313_),
    .Z(_4314_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _4734_ (.A1(_4312_),
    .A2(_4314_),
    .Z(_4315_));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _4735_ (.I(\as2650.carry ),
    .ZN(_4316_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4736_ (.A1(\as2650.psl[3] ),
    .A2(_4316_),
    .ZN(_4317_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _4737_ (.A1(_4317_),
    .A2(_4311_),
    .Z(_4318_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4738_ (.A1(_4315_),
    .A2(_4318_),
    .ZN(_4319_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4739_ (.I(\as2650.psl[3] ),
    .Z(_4320_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4740_ (.A1(_4320_),
    .A2(\as2650.carry ),
    .ZN(_4321_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4741_ (.A1(_4321_),
    .A2(_4311_),
    .ZN(_4322_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4742_ (.I(_4160_),
    .ZN(_4323_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4743_ (.A1(_4323_),
    .A2(_4178_),
    .ZN(_4324_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4744_ (.A1(_4192_),
    .A2(_4324_),
    .ZN(_4325_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_2 _4745_ (.A1(_4303_),
    .A2(_4310_),
    .B(\as2650.psl[3] ),
    .C(\as2650.carry ),
    .ZN(_4326_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _4746_ (.A1(_4322_),
    .A2(_4325_),
    .A3(_4326_),
    .ZN(_4327_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4747_ (.I(_4178_),
    .Z(_4328_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4748_ (.A1(_4323_),
    .A2(_4328_),
    .ZN(_4329_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4749_ (.I(_4329_),
    .Z(_4330_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4750_ (.I(_4257_),
    .Z(_4331_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4751_ (.I(_4331_),
    .Z(_4332_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _4752_ (.I(_4304_),
    .Z(_4333_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4753_ (.I(_4333_),
    .Z(_4334_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _4754_ (.A1(_4332_),
    .A2(_4334_),
    .B(_4309_),
    .ZN(_4335_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4755_ (.I(_4324_),
    .Z(_4336_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _4756_ (.A1(_4290_),
    .A2(_4293_),
    .Z(_4337_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4757_ (.I(_4226_),
    .Z(_4338_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _4758_ (.A1(_4330_),
    .A2(_4335_),
    .B1(_4336_),
    .B2(_4337_),
    .C(_4338_),
    .ZN(_4339_));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _4759_ (.A1(_4319_),
    .A2(_4327_),
    .A3(_4339_),
    .Z(_4340_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _4760_ (.A1(_4183_),
    .A2(_4225_),
    .Z(_4341_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4761_ (.A1(_4341_),
    .A2(_4308_),
    .B(_4279_),
    .ZN(_4342_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _4762_ (.A1(_4279_),
    .A2(_4311_),
    .B1(_4340_),
    .B2(_4342_),
    .ZN(_4343_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4763_ (.I(_4343_),
    .Z(_4344_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4764_ (.I(_4247_),
    .Z(_4345_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4765_ (.I(_4345_),
    .Z(_4346_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4766_ (.I(\as2650.idx_ctrl[0] ),
    .ZN(_4347_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4767_ (.A1(_4243_),
    .A2(_4347_),
    .ZN(_4348_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4768_ (.I(\as2650.idx_ctrl[1] ),
    .ZN(_4349_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4769_ (.A1(_4349_),
    .A2(_4244_),
    .ZN(_4350_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4770_ (.A1(_4348_),
    .A2(_4350_),
    .ZN(_4351_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _4771_ (.A1(_4304_),
    .A2(_4351_),
    .Z(_4352_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4772_ (.I(_4352_),
    .ZN(_4353_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4773_ (.I(_4269_),
    .Z(_4354_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4774_ (.I(\as2650.addr_buff[5] ),
    .ZN(_4355_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4775_ (.A1(\as2650.addr_buff[6] ),
    .A2(_4355_),
    .ZN(_4356_));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _4776_ (.I(\as2650.addr_buff[6] ),
    .ZN(_4357_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _4777_ (.A1(_4357_),
    .A2(\as2650.addr_buff[5] ),
    .ZN(_4358_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _4778_ (.A1(_4356_),
    .A2(_4358_),
    .ZN(_4359_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _4779_ (.A1(_4333_),
    .A2(_4359_),
    .Z(_4360_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4780_ (.I(_4360_),
    .Z(_4361_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4781_ (.I(_4213_),
    .Z(_4362_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4782_ (.I(_4362_),
    .Z(_4363_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4783_ (.I(_4221_),
    .Z(_4364_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4784_ (.I(_4320_),
    .Z(_4365_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4785_ (.I(\as2650.r0[7] ),
    .Z(_4366_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4786_ (.I(_4366_),
    .Z(_4367_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4787_ (.A1(_4367_),
    .A2(_4142_),
    .ZN(_4368_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4788_ (.I(_4298_),
    .Z(_4369_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _4789_ (.I0(\as2650.r123[2][7] ),
    .I1(\as2650.r123_2[2][7] ),
    .S(_4148_),
    .Z(_4370_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4790_ (.A1(_4369_),
    .A2(_4370_),
    .ZN(_4371_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _4791_ (.I0(\as2650.r123[1][7] ),
    .I1(\as2650.r123[0][7] ),
    .I2(\as2650.r123_2[1][7] ),
    .I3(\as2650.r123_2[0][7] ),
    .S0(_4197_),
    .S1(_4148_),
    .Z(_4372_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4792_ (.A1(_4300_),
    .A2(_4372_),
    .ZN(_4373_));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _4793_ (.A1(_4368_),
    .A2(_4371_),
    .A3(_4373_),
    .Z(_4374_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4794_ (.I(_4374_),
    .Z(_4375_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4795_ (.I(_4375_),
    .Z(_4376_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4796_ (.A1(_4365_),
    .A2(_4376_),
    .B(_4321_),
    .ZN(_4377_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4797_ (.I(_4230_),
    .Z(_4378_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4798_ (.I(_4145_),
    .Z(_4379_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _4799_ (.I0(\as2650.r123[2][1] ),
    .I1(\as2650.r123_2[2][1] ),
    .S(_4379_),
    .Z(_4380_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4800_ (.A1(_4297_),
    .A2(_4380_),
    .ZN(_4381_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4801_ (.I(\as2650.r0[1] ),
    .Z(_4382_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4802_ (.I(_4382_),
    .Z(_4383_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _4803_ (.I0(\as2650.r123[1][1] ),
    .I1(\as2650.r123[0][1] ),
    .I2(\as2650.r123_2[1][1] ),
    .I3(\as2650.r123_2[0][1] ),
    .S0(_4139_),
    .S1(_4379_),
    .Z(_4384_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_2 _4804_ (.A1(_4383_),
    .A2(_4140_),
    .B1(_4286_),
    .B2(_4384_),
    .ZN(_4385_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _4805_ (.A1(_4381_),
    .A2(_4385_),
    .Z(_4386_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4806_ (.I(_4386_),
    .Z(_4387_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4807_ (.I(_4387_),
    .Z(_4388_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4808_ (.I(_4229_),
    .Z(_4389_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4809_ (.I(net6),
    .Z(_4390_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4810_ (.I(_4390_),
    .Z(_4391_));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _4811_ (.I(_4391_),
    .ZN(_4392_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _4812_ (.A1(_4172_),
    .A2(_4166_),
    .A3(_4175_),
    .ZN(_4393_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4813_ (.I(_4186_),
    .Z(_4394_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_2 _4814_ (.A1(_4162_),
    .A2(_4393_),
    .A3(_4394_),
    .ZN(_4395_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4815_ (.A1(_4154_),
    .A2(_4395_),
    .ZN(_4396_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4816_ (.I(_4396_),
    .Z(_4397_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _4817_ (.A1(_4216_),
    .A2(_4333_),
    .Z(_4398_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4818_ (.I(_4396_),
    .Z(_4399_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4819_ (.A1(_4398_),
    .A2(_4399_),
    .ZN(_4400_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4820_ (.A1(_4392_),
    .A2(_4397_),
    .B(_4400_),
    .ZN(_4401_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4821_ (.A1(_4389_),
    .A2(_4401_),
    .ZN(_4402_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _4822_ (.A1(_4378_),
    .A2(_4388_),
    .B(_4402_),
    .C(_4222_),
    .ZN(_4403_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4823_ (.A1(_4364_),
    .A2(_4377_),
    .B(_4403_),
    .ZN(_4404_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4824_ (.I(_4285_),
    .Z(_4405_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4825_ (.I(_4405_),
    .Z(_4406_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4826_ (.A1(_4157_),
    .A2(_4268_),
    .ZN(_4407_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4827_ (.A1(_4154_),
    .A2(_4407_),
    .ZN(_4408_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4828_ (.A1(_4406_),
    .A2(_4362_),
    .B(_4408_),
    .ZN(_4409_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _4829_ (.A1(_4363_),
    .A2(_4404_),
    .B(_4409_),
    .ZN(_4410_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _4830_ (.A1(_4354_),
    .A2(_4361_),
    .B(_4410_),
    .C(_4345_),
    .ZN(_4411_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4831_ (.I(_4262_),
    .Z(_4412_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _4832_ (.A1(_4346_),
    .A2(_4353_),
    .B(_4411_),
    .C(_4412_),
    .ZN(_4413_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _4833_ (.A1(_4276_),
    .A2(_4344_),
    .B(_4413_),
    .ZN(_4414_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4834_ (.I(_4205_),
    .Z(_4415_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4835_ (.I(_4415_),
    .Z(_4416_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4836_ (.I(_4170_),
    .Z(_4417_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4837_ (.I(_4417_),
    .Z(_4418_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4838_ (.I(_4418_),
    .Z(_4419_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _4839_ (.I(_4143_),
    .Z(_4420_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4840_ (.I(_4190_),
    .Z(_4421_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _4841_ (.I(_4421_),
    .Z(_4422_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4842_ (.A1(_4224_),
    .A2(_4278_),
    .ZN(_4423_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4843_ (.A1(_4312_),
    .A2(_4423_),
    .ZN(_4424_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4844_ (.I(_4424_),
    .Z(_4425_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _4845_ (.A1(_4420_),
    .A2(_4422_),
    .A3(_4425_),
    .ZN(_4426_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4846_ (.I(_4421_),
    .Z(_4427_));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _4847_ (.I(_4197_),
    .ZN(_4428_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4848_ (.A1(_4428_),
    .A2(_4136_),
    .ZN(_4429_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4849_ (.I(_4429_),
    .Z(_4430_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _4850_ (.A1(_4156_),
    .A2(_4313_),
    .ZN(_4431_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _4851_ (.A1(_4312_),
    .A2(_4431_),
    .ZN(_4432_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _4852_ (.A1(_4427_),
    .A2(_4430_),
    .A3(_4432_),
    .ZN(_4433_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4853_ (.A1(_4426_),
    .A2(_4433_),
    .ZN(_4434_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4854_ (.I(_4434_),
    .Z(_4435_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4855_ (.A1(_4419_),
    .A2(_4435_),
    .ZN(_4436_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4856_ (.I(_4436_),
    .ZN(_4437_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4857_ (.I(_4202_),
    .Z(_4438_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_2 _4858_ (.A1(_4416_),
    .A2(_4437_),
    .B(_4273_),
    .C(_4438_),
    .ZN(_4439_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4859_ (.I(_4439_),
    .Z(_4440_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4860_ (.I(_4406_),
    .Z(_4441_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4861_ (.I(_4211_),
    .Z(_4442_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4862_ (.I(_4442_),
    .Z(_4443_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _4863_ (.A1(_4443_),
    .A2(_4426_),
    .ZN(_4444_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4864_ (.A1(_4415_),
    .A2(_4444_),
    .ZN(_4445_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4865_ (.I(_4445_),
    .ZN(_4446_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4866_ (.A1(_4441_),
    .A2(_4446_),
    .ZN(_4447_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4867_ (.I(\as2650.psu[2] ),
    .Z(_4448_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4868_ (.A1(\as2650.psu[0] ),
    .A2(\as2650.psu[1] ),
    .ZN(_4449_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4869_ (.I(_4449_),
    .Z(_4450_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4870_ (.A1(_4448_),
    .A2(_4450_),
    .ZN(_4451_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4871_ (.I(_4451_),
    .Z(_4452_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _4872_ (.A1(\as2650.psu[2] ),
    .A2(_4449_),
    .Z(_4453_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4873_ (.I(_4453_),
    .Z(_4454_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4874_ (.A1(\as2650.stack[3][8] ),
    .A2(_4452_),
    .B(_4454_),
    .ZN(_4455_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4875_ (.I(\as2650.psu[0] ),
    .ZN(_4456_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4876_ (.I(\as2650.psu[1] ),
    .ZN(_4457_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4877_ (.I(_4457_),
    .Z(_4458_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4878_ (.A1(_4456_),
    .A2(_4458_),
    .ZN(_4459_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4879_ (.I(_4459_),
    .Z(_4460_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4880_ (.I(_4460_),
    .Z(_4461_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4881_ (.A1(\as2650.stack[2][8] ),
    .A2(_4461_),
    .ZN(_4462_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4882_ (.I(\as2650.psu[1] ),
    .Z(_4463_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4883_ (.A1(_4456_),
    .A2(_4463_),
    .ZN(_4464_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4884_ (.I(_4464_),
    .Z(_4465_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4885_ (.I(_4465_),
    .Z(_4466_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4886_ (.I(\as2650.psu[0] ),
    .Z(_4467_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4887_ (.A1(_4467_),
    .A2(_4458_),
    .ZN(_4468_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4888_ (.I(_4468_),
    .Z(_4469_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4889_ (.I(_4469_),
    .Z(_4470_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _4890_ (.A1(\as2650.stack[0][8] ),
    .A2(_4466_),
    .B1(_4470_),
    .B2(\as2650.stack[1][8] ),
    .ZN(_4471_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _4891_ (.A1(_4455_),
    .A2(_4462_),
    .A3(_4471_),
    .ZN(_4472_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4892_ (.A1(_4448_),
    .A2(_4450_),
    .ZN(_4473_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _4893_ (.A1(_4448_),
    .A2(_4449_),
    .Z(_4474_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4894_ (.A1(_4473_),
    .A2(_4474_),
    .ZN(_4475_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4895_ (.I(_4475_),
    .Z(_4476_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4896_ (.I(_4476_),
    .Z(_4477_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4897_ (.I(_4450_),
    .Z(_4478_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4898_ (.I(_4478_),
    .Z(_4479_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _4899_ (.A1(\as2650.stack[7][8] ),
    .A2(_4479_),
    .B1(_4461_),
    .B2(\as2650.stack[6][8] ),
    .ZN(_4480_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4900_ (.I(_4464_),
    .Z(_4481_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4901_ (.I(_4481_),
    .Z(_4482_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _4902_ (.A1(\as2650.stack[4][8] ),
    .A2(_4482_),
    .B1(_4470_),
    .B2(\as2650.stack[5][8] ),
    .ZN(_4483_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _4903_ (.A1(_4477_),
    .A2(_4480_),
    .A3(_4483_),
    .ZN(_4484_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4904_ (.I(_4445_),
    .Z(_4485_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _4905_ (.A1(_4472_),
    .A2(_4484_),
    .B(_4485_),
    .ZN(_4486_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4906_ (.I(_4211_),
    .Z(_4487_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4907_ (.I(_4191_),
    .Z(_4488_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _4908_ (.A1(_4143_),
    .A2(_4488_),
    .A3(_4432_),
    .ZN(_4489_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _4909_ (.A1(_4487_),
    .A2(_4489_),
    .Z(_4490_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4910_ (.I(_4490_),
    .Z(_4491_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4911_ (.A1(_4436_),
    .A2(_4491_),
    .ZN(_4492_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4912_ (.A1(_4415_),
    .A2(_4492_),
    .ZN(_4493_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4913_ (.I(_4493_),
    .Z(_4494_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_1 _4914_ (.A1(_4439_),
    .A2(_4447_),
    .A3(_4486_),
    .A4(_4494_),
    .ZN(_4495_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _4915_ (.A1(\as2650.r123[0][0] ),
    .A2(_4440_),
    .B(_4495_),
    .ZN(_4496_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4916_ (.A1(_4275_),
    .A2(_4414_),
    .B(_4496_),
    .ZN(_0000_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4917_ (.I(\as2650.r123[0][1] ),
    .ZN(_4497_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4918_ (.I(_4439_),
    .Z(_4498_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4919_ (.I(_4498_),
    .Z(_4499_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4920_ (.I(_4274_),
    .Z(_4500_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4921_ (.I(_4408_),
    .Z(_4501_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4922_ (.I(_4356_),
    .Z(_4502_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _4923_ (.A1(\as2650.addr_buff[6] ),
    .A2(_4355_),
    .ZN(_4503_));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _4924_ (.A1(_4305_),
    .A2(_4306_),
    .A3(_4503_),
    .Z(_4504_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_2 _4925_ (.A1(_4283_),
    .A2(_4289_),
    .B1(_4381_),
    .B2(_4385_),
    .ZN(_4505_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4926_ (.I(_4505_),
    .Z(_4506_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4927_ (.I(_4506_),
    .Z(_4507_));
 gf180mcu_fd_sc_mcu7t5v0__and4_1 _4928_ (.A1(_4282_),
    .A2(_4288_),
    .A3(_4381_),
    .A4(_4385_),
    .Z(_4508_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4929_ (.I(_4508_),
    .Z(_4509_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4930_ (.I(_4509_),
    .Z(_4510_));
 gf180mcu_fd_sc_mcu7t5v0__or4_1 _4931_ (.A1(_4502_),
    .A2(_4504_),
    .A3(_4507_),
    .A4(_4510_),
    .Z(_4511_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _4932_ (.A1(_4502_),
    .A2(_4504_),
    .B1(_4507_),
    .B2(_4510_),
    .ZN(_4512_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _4933_ (.A1(_4511_),
    .A2(_4512_),
    .Z(_4513_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4934_ (.A1(_4305_),
    .A2(_4306_),
    .ZN(_4514_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4935_ (.I(_4389_),
    .Z(_4515_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _4936_ (.I(_4147_),
    .Z(_4516_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _4937_ (.I0(\as2650.r123[2][2] ),
    .I1(\as2650.r123_2[2][2] ),
    .S(_4516_),
    .Z(_4517_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4938_ (.A1(_4297_),
    .A2(_4517_),
    .ZN(_4518_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4939_ (.I(\as2650.r0[2] ),
    .Z(_4519_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4940_ (.I(_4519_),
    .Z(_4520_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4941_ (.I(_4286_),
    .Z(_4521_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_2 _4942_ (.I0(\as2650.r123[1][2] ),
    .I1(\as2650.r123[0][2] ),
    .I2(\as2650.r123_2[1][2] ),
    .I3(\as2650.r123_2[0][2] ),
    .S0(_4139_),
    .S1(_4379_),
    .Z(_4522_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_2 _4943_ (.A1(_4520_),
    .A2(_4140_),
    .B1(_4521_),
    .B2(_4522_),
    .ZN(_4523_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _4944_ (.A1(_4518_),
    .A2(_4523_),
    .Z(_4524_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4945_ (.I(_4524_),
    .Z(_4525_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4946_ (.I(_4525_),
    .Z(_4526_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4947_ (.I(_4526_),
    .Z(_4527_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4948_ (.I(net7),
    .Z(_4528_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4949_ (.I(_4528_),
    .Z(_4529_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4950_ (.I(_4529_),
    .Z(_4530_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4951_ (.I(_4530_),
    .Z(_4531_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4952_ (.I(_4399_),
    .Z(_4532_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _4953_ (.A1(_4249_),
    .A2(_4258_),
    .ZN(_4533_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _4954_ (.I0(_4217_),
    .I1(_4533_),
    .S(_4333_),
    .Z(_4534_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _4955_ (.A1(_4387_),
    .A2(_4534_),
    .Z(_4535_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4956_ (.A1(_4397_),
    .A2(_4535_),
    .ZN(_4536_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _4957_ (.A1(_4531_),
    .A2(_4532_),
    .B(_4536_),
    .C(_4231_),
    .ZN(_4537_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4958_ (.I(_4221_),
    .Z(_4538_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _4959_ (.A1(_4515_),
    .A2(_4527_),
    .B(_4537_),
    .C(_4538_),
    .ZN(_4539_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _4960_ (.A1(_4364_),
    .A2(_4514_),
    .B(_4539_),
    .C(_4363_),
    .ZN(_4540_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4961_ (.I(_4383_),
    .Z(_4541_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4962_ (.I(_4541_),
    .Z(_4542_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _4963_ (.I(_4487_),
    .Z(_4543_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _4964_ (.A1(_4422_),
    .A2(_4194_),
    .ZN(_4544_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_2 _4965_ (.A1(_4206_),
    .A2(_4543_),
    .A3(_4544_),
    .ZN(_4545_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4966_ (.I(_4545_),
    .Z(_4546_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4967_ (.I(_4546_),
    .Z(_4547_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4968_ (.A1(_4542_),
    .A2(_4547_),
    .ZN(_4548_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _4969_ (.A1(_4501_),
    .A2(_4540_),
    .A3(_4548_),
    .ZN(_4549_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4970_ (.I(_4232_),
    .Z(_4550_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _4971_ (.I(_4550_),
    .Z(_4551_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _4972_ (.A1(_4551_),
    .A2(_4242_),
    .A3(_4246_),
    .ZN(_4552_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4973_ (.A1(_4154_),
    .A2(_4552_),
    .ZN(_0284_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4974_ (.I(_0284_),
    .Z(_0285_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _4975_ (.A1(_4501_),
    .A2(_4513_),
    .B(_4549_),
    .C(_0285_),
    .ZN(_0286_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4976_ (.A1(_4243_),
    .A2(_4347_),
    .ZN(_0287_));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _4977_ (.A1(_4305_),
    .A2(_4306_),
    .A3(_0287_),
    .Z(_0288_));
 gf180mcu_fd_sc_mcu7t5v0__or4_1 _4978_ (.A1(_4348_),
    .A2(_0288_),
    .A3(_4506_),
    .A4(_4509_),
    .Z(_0289_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4979_ (.I(_4508_),
    .Z(_0290_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _4980_ (.A1(_4348_),
    .A2(_0288_),
    .B1(_4506_),
    .B2(_0290_),
    .ZN(_0291_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _4981_ (.A1(_0289_),
    .A2(_0291_),
    .Z(_0292_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _4982_ (.A1(_4346_),
    .A2(_0292_),
    .B(_4412_),
    .ZN(_0293_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4983_ (.I(_4248_),
    .Z(_0294_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _4984_ (.A1(_0294_),
    .A2(_4261_),
    .Z(_0295_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4985_ (.I(_0295_),
    .Z(_0296_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4986_ (.I(\as2650.holding_reg[1] ),
    .Z(_0297_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4987_ (.A1(_4257_),
    .A2(_4386_),
    .ZN(_0298_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4988_ (.A1(_0297_),
    .A2(_4332_),
    .B(_0298_),
    .ZN(_0299_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4989_ (.A1(_4279_),
    .A2(_0299_),
    .ZN(_0300_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4990_ (.A1(_4381_),
    .A2(_4385_),
    .ZN(_0301_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4991_ (.A1(\as2650.holding_reg[1] ),
    .A2(_0301_),
    .ZN(_0302_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4992_ (.I(_0302_),
    .Z(_0303_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _4993_ (.A1(\as2650.holding_reg[1] ),
    .A2(_0301_),
    .Z(_0304_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4994_ (.A1(_0302_),
    .A2(_0304_),
    .ZN(_0305_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _4995_ (.A1(_4290_),
    .A2(_4293_),
    .A3(_4302_),
    .ZN(_0306_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _4996_ (.A1(_4317_),
    .A2(_0306_),
    .B(_4310_),
    .ZN(_0307_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _4997_ (.A1(_0305_),
    .A2(_0307_),
    .Z(_0308_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4998_ (.A1(_4315_),
    .A2(_0308_),
    .ZN(_0309_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _4999_ (.A1(_4302_),
    .A2(_4326_),
    .B(_0305_),
    .ZN(_0310_));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _5000_ (.A1(_4302_),
    .A2(_4326_),
    .A3(_0305_),
    .Z(_0311_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5001_ (.A1(_0310_),
    .A2(_0311_),
    .B(_4325_),
    .ZN(_0312_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5002_ (.A1(_4277_),
    .A2(_4329_),
    .ZN(_0313_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5003_ (.I(_4331_),
    .Z(_0314_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5004_ (.A1(_0297_),
    .A2(_0314_),
    .ZN(_0315_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _5005_ (.A1(_4332_),
    .A2(_4386_),
    .B(_4324_),
    .C(_0315_),
    .ZN(_0316_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _5006_ (.A1(_0309_),
    .A2(_0312_),
    .A3(_0313_),
    .A4(_0316_),
    .ZN(_0317_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _5007_ (.A1(_4330_),
    .A2(_0304_),
    .B(_4338_),
    .ZN(_0318_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _5008_ (.A1(_4338_),
    .A2(_0303_),
    .B1(_0317_),
    .B2(_0318_),
    .ZN(_0319_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _5009_ (.A1(_0300_),
    .A2(_0319_),
    .Z(_0320_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5010_ (.I(_0320_),
    .Z(_0321_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5011_ (.A1(_0296_),
    .A2(_0321_),
    .ZN(_0322_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _5012_ (.A1(_0286_),
    .A2(_0293_),
    .B(_0322_),
    .ZN(_0323_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5013_ (.I(_4468_),
    .Z(_0324_));
 gf180mcu_fd_sc_mcu7t5v0__aoi222_2 _5014_ (.A1(\as2650.stack[4][9] ),
    .A2(_4481_),
    .B1(_4460_),
    .B2(\as2650.stack[6][9] ),
    .C1(_0324_),
    .C2(\as2650.stack[5][9] ),
    .ZN(_0325_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5015_ (.I(_4478_),
    .Z(_0326_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5016_ (.A1(_4453_),
    .A2(_4451_),
    .ZN(_0327_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5017_ (.I(_0327_),
    .Z(_0328_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5018_ (.I(_0328_),
    .Z(_0329_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _5019_ (.A1(\as2650.stack[7][9] ),
    .A2(_0326_),
    .B(_0329_),
    .ZN(_0330_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5020_ (.A1(\as2650.stack[3][9] ),
    .A2(_4452_),
    .B(_4454_),
    .ZN(_0331_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5021_ (.A1(\as2650.stack[2][9] ),
    .A2(_4460_),
    .ZN(_0332_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _5022_ (.A1(\as2650.stack[0][9] ),
    .A2(_4465_),
    .B1(_0324_),
    .B2(\as2650.stack[1][9] ),
    .ZN(_0333_));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _5023_ (.A1(_0331_),
    .A2(_0332_),
    .A3(_0333_),
    .Z(_0334_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _5024_ (.A1(_0325_),
    .A2(_0330_),
    .B(_0334_),
    .ZN(_0335_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5025_ (.A1(_4485_),
    .A2(_0335_),
    .ZN(_0336_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5026_ (.I(_4542_),
    .Z(_0337_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5027_ (.A1(_4420_),
    .A2(_4488_),
    .ZN(_0338_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _5028_ (.I(_0338_),
    .Z(_0339_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _5029_ (.A1(_4277_),
    .A2(_4423_),
    .Z(_0340_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5030_ (.A1(_0339_),
    .A2(_0340_),
    .ZN(_0341_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5031_ (.I(_0341_),
    .Z(_0342_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5032_ (.I(_0342_),
    .Z(_0343_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5033_ (.A1(_0337_),
    .A2(_0343_),
    .ZN(_0344_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _5034_ (.A1(_4494_),
    .A2(_0336_),
    .A3(_0344_),
    .ZN(_0345_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _5035_ (.A1(_4500_),
    .A2(_0323_),
    .B(_0345_),
    .C(_4498_),
    .ZN(_0346_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _5036_ (.A1(_4497_),
    .A2(_4499_),
    .B(_0346_),
    .ZN(_0001_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5037_ (.I(\as2650.r123[0][2] ),
    .ZN(_0347_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5038_ (.I(_0287_),
    .Z(_0348_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5039_ (.A1(_4518_),
    .A2(_4523_),
    .ZN(_0349_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_2 _5040_ (.A1(_0349_),
    .A2(_4509_),
    .Z(_0350_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _5041_ (.A1(_0348_),
    .A2(_0350_),
    .ZN(_0351_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _5042_ (.A1(_4349_),
    .A2(_4244_),
    .ZN(_0352_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5043_ (.A1(_0352_),
    .A2(_0287_),
    .ZN(_0353_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5044_ (.I(_0349_),
    .Z(_0354_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _5045_ (.I(_0354_),
    .Z(_0355_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_2 _5046_ (.A1(_0349_),
    .A2(_4505_),
    .Z(_0356_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_4 _5047_ (.A1(_0353_),
    .A2(_0355_),
    .B1(_0356_),
    .B2(_0352_),
    .ZN(_0357_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _5048_ (.A1(_0351_),
    .A2(_0357_),
    .ZN(_0358_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5049_ (.I(_4520_),
    .Z(_0359_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5050_ (.I(_0359_),
    .Z(_0360_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5051_ (.I(_0360_),
    .Z(_0361_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5052_ (.I(\as2650.r0[3] ),
    .Z(_0362_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5053_ (.I(_0362_),
    .Z(_0363_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5054_ (.I(_0363_),
    .Z(_0364_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5055_ (.A1(_0364_),
    .A2(_4141_),
    .ZN(_0365_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _5056_ (.I0(\as2650.r123[2][3] ),
    .I1(\as2650.r123_2[2][3] ),
    .S(_4516_),
    .Z(_0366_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _5057_ (.I0(\as2650.r123[1][3] ),
    .I1(\as2650.r123[0][3] ),
    .I2(\as2650.r123_2[1][3] ),
    .I3(\as2650.r123_2[0][3] ),
    .S0(_4139_),
    .S1(_4516_),
    .Z(_0367_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _5058_ (.A1(_4297_),
    .A2(_0366_),
    .B1(_0367_),
    .B2(_4521_),
    .ZN(_0368_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5059_ (.A1(_0365_),
    .A2(_0368_),
    .ZN(_0369_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5060_ (.I(_0369_),
    .Z(_0370_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5061_ (.I(_0370_),
    .Z(_0371_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5062_ (.I(_0371_),
    .Z(_0372_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5063_ (.I(net8),
    .Z(_0373_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _5064_ (.I(_0373_),
    .ZN(_0374_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5065_ (.I(_0374_),
    .Z(_0375_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5066_ (.I(_0375_),
    .Z(_0376_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _5067_ (.A1(_4218_),
    .A2(_4507_),
    .B1(_4510_),
    .B2(_4533_),
    .ZN(_0377_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _5068_ (.A1(_4525_),
    .A2(_0377_),
    .Z(_0378_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5069_ (.A1(_4399_),
    .A2(_0378_),
    .ZN(_0379_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _5070_ (.A1(_0376_),
    .A2(_4397_),
    .B(_0379_),
    .C(_4230_),
    .ZN(_0380_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _5071_ (.A1(_4378_),
    .A2(_0372_),
    .B(_0380_),
    .C(_4222_),
    .ZN(_0381_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _5072_ (.A1(_4538_),
    .A2(_4388_),
    .B(_0381_),
    .C(_4362_),
    .ZN(_0382_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _5073_ (.A1(_0361_),
    .A2(_4363_),
    .B(_4408_),
    .C(_0382_),
    .ZN(_0383_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5074_ (.I(_4503_),
    .Z(_0384_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5075_ (.A1(_0384_),
    .A2(_0350_),
    .ZN(_0385_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5076_ (.A1(_4357_),
    .A2(\as2650.addr_buff[5] ),
    .ZN(_0386_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5077_ (.A1(_4359_),
    .A2(_4525_),
    .ZN(_0387_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5078_ (.A1(_0386_),
    .A2(_0356_),
    .B(_0387_),
    .ZN(_0388_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5079_ (.A1(_0385_),
    .A2(_0388_),
    .ZN(_0389_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5080_ (.A1(_4354_),
    .A2(_0389_),
    .ZN(_0390_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _5081_ (.A1(_0383_),
    .A2(_0390_),
    .B(_4345_),
    .ZN(_0391_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _5082_ (.A1(_4346_),
    .A2(_0358_),
    .B(_0391_),
    .ZN(_0392_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5083_ (.I(_4312_),
    .Z(_0393_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5084_ (.I(_4278_),
    .Z(_0394_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _5085_ (.A1(_0393_),
    .A2(_0394_),
    .Z(_0395_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5086_ (.I(_0395_),
    .Z(_0396_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _5087_ (.I(_4341_),
    .Z(_0397_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _5088_ (.A1(\as2650.holding_reg[2] ),
    .A2(_0355_),
    .Z(_0398_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _5089_ (.A1(\as2650.holding_reg[2] ),
    .A2(_0355_),
    .Z(_0399_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5090_ (.I(_0354_),
    .Z(_0400_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5091_ (.A1(\as2650.holding_reg[2] ),
    .A2(_0400_),
    .ZN(_0401_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _5092_ (.A1(_0401_),
    .A2(_0399_),
    .Z(_0402_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _5093_ (.A1(_0303_),
    .A2(_0304_),
    .Z(_0403_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _5094_ (.A1(_0297_),
    .A2(_4331_),
    .B(_0298_),
    .C(_0303_),
    .ZN(_0404_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5095_ (.A1(_0403_),
    .A2(_0307_),
    .B(_0404_),
    .ZN(_0405_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _5096_ (.A1(_0402_),
    .A2(_0405_),
    .Z(_0406_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5097_ (.I(_0303_),
    .ZN(_0407_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5098_ (.I(_0402_),
    .Z(_0408_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5099_ (.A1(_0407_),
    .A2(_0310_),
    .B(_0408_),
    .ZN(_0409_));
 gf180mcu_fd_sc_mcu7t5v0__or3_1 _5100_ (.A1(_0407_),
    .A2(_0310_),
    .A3(_0408_),
    .Z(_0410_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _5101_ (.A1(_4277_),
    .A2(_4324_),
    .Z(_0411_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _5102_ (.A1(_0409_),
    .A2(_0410_),
    .B(_0411_),
    .ZN(_0412_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5103_ (.I(\as2650.holding_reg[2] ),
    .Z(_0413_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5104_ (.I(_0314_),
    .Z(_0414_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5105_ (.A1(_0414_),
    .A2(_4526_),
    .ZN(_0415_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _5106_ (.A1(_0413_),
    .A2(_0414_),
    .B(_4314_),
    .C(_0415_),
    .ZN(_0416_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _5107_ (.A1(_4315_),
    .A2(_0406_),
    .B(_0412_),
    .C(_0416_),
    .ZN(_0417_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5108_ (.I(_4330_),
    .Z(_0418_));
 gf180mcu_fd_sc_mcu7t5v0__oai222_1 _5109_ (.A1(_0397_),
    .A2(_0398_),
    .B1(_0399_),
    .B2(_0313_),
    .C1(_0417_),
    .C2(_0418_),
    .ZN(_0419_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5110_ (.A1(_0395_),
    .A2(_0408_),
    .ZN(_0420_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5111_ (.A1(_0396_),
    .A2(_0419_),
    .B(_0420_),
    .ZN(_0421_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5112_ (.I(_0421_),
    .Z(_0422_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5113_ (.A1(_4276_),
    .A2(_0422_),
    .ZN(_0423_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _5114_ (.A1(_4276_),
    .A2(_0392_),
    .B(_0423_),
    .ZN(_0424_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5115_ (.A1(\as2650.stack[3][10] ),
    .A2(_4452_),
    .B(_4454_),
    .ZN(_0425_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5116_ (.I(_4459_),
    .Z(_0426_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5117_ (.I(_0426_),
    .Z(_0427_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5118_ (.A1(\as2650.stack[2][10] ),
    .A2(_0427_),
    .ZN(_0428_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5119_ (.I(_4465_),
    .Z(_0429_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5120_ (.I(_4469_),
    .Z(_0430_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _5121_ (.A1(\as2650.stack[0][10] ),
    .A2(_0429_),
    .B1(_0430_),
    .B2(\as2650.stack[1][10] ),
    .ZN(_0431_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _5122_ (.A1(_0425_),
    .A2(_0428_),
    .A3(_0431_),
    .ZN(_0432_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _5123_ (.A1(\as2650.stack[4][10] ),
    .A2(_0429_),
    .B1(_4470_),
    .B2(\as2650.stack[5][10] ),
    .ZN(_0433_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _5124_ (.A1(\as2650.stack[7][10] ),
    .A2(_0326_),
    .B1(_0427_),
    .B2(\as2650.stack[6][10] ),
    .ZN(_0434_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _5125_ (.A1(_4477_),
    .A2(_0433_),
    .A3(_0434_),
    .ZN(_0435_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5126_ (.A1(_0432_),
    .A2(_0435_),
    .ZN(_0436_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5127_ (.A1(_0361_),
    .A2(_0342_),
    .ZN(_0437_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5128_ (.I(_4493_),
    .Z(_0438_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _5129_ (.A1(_4446_),
    .A2(_0436_),
    .B(_0437_),
    .C(_0438_),
    .ZN(_0439_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _5130_ (.A1(_4500_),
    .A2(_0424_),
    .B(_0439_),
    .C(_4498_),
    .ZN(_0440_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _5131_ (.A1(_0347_),
    .A2(_4499_),
    .B(_0440_),
    .ZN(_0002_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5132_ (.I(\as2650.r123[0][3] ),
    .ZN(_0441_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _5133_ (.A1(\as2650.holding_reg[3] ),
    .A2(_0370_),
    .Z(_0442_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5134_ (.A1(\as2650.holding_reg[3] ),
    .A2(_0371_),
    .ZN(_0443_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5135_ (.A1(_0442_),
    .A2(_0443_),
    .ZN(_0444_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5136_ (.I(_0444_),
    .Z(_0445_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5137_ (.A1(_0395_),
    .A2(_0445_),
    .ZN(_0446_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5138_ (.I(_0393_),
    .Z(_0447_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5139_ (.A1(_0447_),
    .A2(_4314_),
    .ZN(_0448_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5140_ (.A1(_0401_),
    .A2(_0399_),
    .ZN(_0449_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5141_ (.A1(_4257_),
    .A2(_4525_),
    .ZN(_0450_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5142_ (.A1(_0413_),
    .A2(_4331_),
    .B(_0450_),
    .ZN(_0451_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5143_ (.A1(_0398_),
    .A2(_0451_),
    .ZN(_0452_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _5144_ (.A1(_0449_),
    .A2(_0405_),
    .B(_0452_),
    .ZN(_0453_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _5145_ (.A1(_0445_),
    .A2(_0453_),
    .ZN(_0454_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5146_ (.A1(_0448_),
    .A2(_0454_),
    .ZN(_0455_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _5147_ (.A1(_4300_),
    .A2(_4522_),
    .Z(_0456_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5148_ (.A1(_0359_),
    .A2(_4142_),
    .ZN(_0457_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5149_ (.A1(_4518_),
    .A2(_0457_),
    .ZN(_0458_));
 gf180mcu_fd_sc_mcu7t5v0__oai33_1 _5150_ (.A1(_0413_),
    .A2(_0456_),
    .A3(_0458_),
    .B1(_0407_),
    .B2(_0310_),
    .B3(_0398_),
    .ZN(_0459_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _5151_ (.A1(_0444_),
    .A2(_0459_),
    .Z(_0460_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5152_ (.I(\as2650.holding_reg[3] ),
    .Z(_0461_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _5153_ (.A1(_0365_),
    .A2(_0368_),
    .Z(_0462_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5154_ (.I(_0462_),
    .Z(_0463_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _5155_ (.I(_0463_),
    .Z(_0464_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5156_ (.A1(_0314_),
    .A2(_0464_),
    .ZN(_0465_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5157_ (.A1(_0461_),
    .A2(_0314_),
    .B(_0465_),
    .ZN(_0466_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5158_ (.I(_0466_),
    .Z(_0467_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _5159_ (.A1(_0393_),
    .A2(_0467_),
    .Z(_0468_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5160_ (.I(_4191_),
    .Z(_0469_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5161_ (.A1(_0469_),
    .A2(_0464_),
    .ZN(_0470_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _5162_ (.A1(_0461_),
    .A2(_4422_),
    .B(_4336_),
    .C(_0470_),
    .ZN(_0471_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_2 _5163_ (.A1(_0411_),
    .A2(_0460_),
    .B1(_0468_),
    .B2(_4225_),
    .C(_0471_),
    .ZN(_0472_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _5164_ (.I(_4279_),
    .Z(_0473_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_2 _5165_ (.A1(_0397_),
    .A2(_0442_),
    .B1(_0455_),
    .B2(_0472_),
    .C(_0473_),
    .ZN(_0474_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5166_ (.A1(_0446_),
    .A2(_0474_),
    .ZN(_0475_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5167_ (.I(_0475_),
    .Z(_0476_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _5168_ (.A1(_0354_),
    .A2(_4505_),
    .A3(_0369_),
    .ZN(_0477_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_1 _5169_ (.A1(_4304_),
    .A2(_4386_),
    .A3(_4524_),
    .B(_0463_),
    .ZN(_0478_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _5170_ (.A1(_0477_),
    .A2(_0478_),
    .B(_0352_),
    .ZN(_0479_));
 gf180mcu_fd_sc_mcu7t5v0__and4_1 _5171_ (.A1(_4518_),
    .A2(_4523_),
    .A3(_0365_),
    .A4(_0368_),
    .Z(_0480_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5172_ (.I(_0480_),
    .Z(_0481_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _5173_ (.A1(_4509_),
    .A2(_0481_),
    .Z(_0482_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _5174_ (.A1(_4524_),
    .A2(_0290_),
    .B(_0462_),
    .ZN(_0483_));
 gf180mcu_fd_sc_mcu7t5v0__oai32_1 _5175_ (.A1(_0348_),
    .A2(_0482_),
    .A3(_0483_),
    .B1(_0353_),
    .B2(_0370_),
    .ZN(_0484_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _5176_ (.A1(_0479_),
    .A2(_0484_),
    .Z(_0485_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5177_ (.I(_4269_),
    .Z(_0486_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _5178_ (.I(_4359_),
    .Z(_0487_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5179_ (.A1(_0477_),
    .A2(_0478_),
    .ZN(_0488_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_2 _5180_ (.A1(_0384_),
    .A2(_0482_),
    .A3(_0483_),
    .ZN(_0489_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_4 _5181_ (.A1(_0487_),
    .A2(_0464_),
    .B1(_0488_),
    .B2(_4502_),
    .C(_0489_),
    .ZN(_0490_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5182_ (.I(_0490_),
    .Z(_0491_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5183_ (.I(_0364_),
    .Z(_0492_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _5184_ (.I(_4379_),
    .Z(_0493_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _5185_ (.I0(\as2650.r123[1][4] ),
    .I1(\as2650.r123[0][4] ),
    .I2(\as2650.r123_2[1][4] ),
    .I3(\as2650.r123_2[0][4] ),
    .S0(_4196_),
    .S1(_0493_),
    .Z(_0494_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5186_ (.A1(_4521_),
    .A2(_0494_),
    .ZN(_0495_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _5187_ (.I0(\as2650.r123[2][4] ),
    .I1(\as2650.r123_2[2][4] ),
    .S(_4516_),
    .Z(_0496_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5188_ (.A1(_4298_),
    .A2(_0496_),
    .ZN(_0497_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5189_ (.I(\as2650.r0[4] ),
    .Z(_0498_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5190_ (.I(_0498_),
    .Z(_0499_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5191_ (.I(_0499_),
    .Z(_0500_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5192_ (.A1(_0500_),
    .A2(_4141_),
    .ZN(_0501_));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _5193_ (.A1(_0495_),
    .A2(_0497_),
    .A3(_0501_),
    .Z(_0502_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5194_ (.I(_0502_),
    .Z(_0503_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5195_ (.I(_0503_),
    .Z(_0504_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5196_ (.I(_0504_),
    .Z(_0505_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5197_ (.I(net9),
    .Z(_0506_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5198_ (.I(_0506_),
    .Z(_0507_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5199_ (.I(_0507_),
    .Z(_0508_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _5200_ (.A1(_4218_),
    .A2(_0355_),
    .A3(_4507_),
    .ZN(_0509_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _5201_ (.A1(_4533_),
    .A2(_4524_),
    .A3(_4510_),
    .ZN(_0510_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5202_ (.A1(_0509_),
    .A2(_0510_),
    .ZN(_0511_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_2 _5203_ (.A1(_0463_),
    .A2(_0511_),
    .Z(_0512_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5204_ (.A1(_4396_),
    .A2(_0512_),
    .ZN(_0513_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _5205_ (.A1(_0508_),
    .A2(_4399_),
    .B(_0513_),
    .C(_4230_),
    .ZN(_0514_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _5206_ (.A1(_4389_),
    .A2(_0505_),
    .B(_0514_),
    .C(_4221_),
    .ZN(_0515_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5207_ (.I(_4220_),
    .Z(_0516_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _5208_ (.A1(_4212_),
    .A2(_0516_),
    .Z(_0517_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _5209_ (.A1(_0517_),
    .A2(_4526_),
    .B(_4545_),
    .ZN(_0518_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _5210_ (.A1(_0492_),
    .A2(_4545_),
    .B1(_0515_),
    .B2(_0518_),
    .ZN(_0519_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5211_ (.A1(_4269_),
    .A2(_0519_),
    .ZN(_0520_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _5212_ (.A1(_0486_),
    .A2(_0491_),
    .B(_0520_),
    .C(_4247_),
    .ZN(_0521_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _5213_ (.A1(_4345_),
    .A2(_0485_),
    .B(_0521_),
    .C(_4262_),
    .ZN(_0522_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _5214_ (.A1(_4412_),
    .A2(_0476_),
    .B(_0522_),
    .ZN(_0523_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5215_ (.I(_0523_),
    .ZN(_0524_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5216_ (.I(_0328_),
    .Z(_0525_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _5217_ (.I(_0525_),
    .Z(_0526_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _5218_ (.I(_0426_),
    .Z(_0527_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _5219_ (.A1(\as2650.stack[3][11] ),
    .A2(_4450_),
    .B1(_4469_),
    .B2(\as2650.stack[1][11] ),
    .ZN(_0528_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5220_ (.I(_0528_),
    .ZN(_0529_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_2 _5221_ (.A1(\as2650.stack[0][11] ),
    .A2(_0429_),
    .B1(_0527_),
    .B2(\as2650.stack[2][11] ),
    .C(_0529_),
    .ZN(_0530_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _5222_ (.A1(\as2650.stack[4][11] ),
    .A2(_0429_),
    .B1(_0430_),
    .B2(\as2650.stack[5][11] ),
    .ZN(_0531_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_2 _5223_ (.A1(\as2650.stack[7][11] ),
    .A2(_4478_),
    .B1(_0527_),
    .B2(\as2650.stack[6][11] ),
    .C(_0329_),
    .ZN(_0532_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_2 _5224_ (.A1(_0526_),
    .A2(_0530_),
    .B1(_0531_),
    .B2(_0532_),
    .ZN(_0533_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5225_ (.A1(_4485_),
    .A2(_0533_),
    .ZN(_0534_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5226_ (.I(_0492_),
    .Z(_0535_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5227_ (.A1(_0535_),
    .A2(_0343_),
    .ZN(_0536_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _5228_ (.A1(_4494_),
    .A2(_0534_),
    .A3(_0536_),
    .ZN(_0537_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5229_ (.I(_4439_),
    .Z(_0538_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _5230_ (.A1(_4500_),
    .A2(_0524_),
    .B(_0537_),
    .C(_0538_),
    .ZN(_0539_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _5231_ (.A1(_0441_),
    .A2(_4499_),
    .B(_0539_),
    .ZN(_0003_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5232_ (.I(\as2650.r123[0][4] ),
    .ZN(_0540_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _5233_ (.A1(_0495_),
    .A2(_0497_),
    .A3(_0501_),
    .ZN(_0541_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5234_ (.I(_0541_),
    .Z(_0542_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _5235_ (.A1(\as2650.holding_reg[4] ),
    .A2(_0542_),
    .Z(_0543_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5236_ (.I(_4325_),
    .Z(_0544_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5237_ (.A1(_0461_),
    .A2(_0371_),
    .ZN(_0545_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5238_ (.A1(_0443_),
    .A2(_0459_),
    .B(_0545_),
    .ZN(_0546_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _5239_ (.A1(_0543_),
    .A2(_0546_),
    .Z(_0547_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5240_ (.I(_0414_),
    .Z(_0548_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5241_ (.I(\as2650.holding_reg[4] ),
    .Z(_0549_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5242_ (.I(_4332_),
    .Z(_0550_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5243_ (.A1(_0549_),
    .A2(_0550_),
    .ZN(_0551_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5244_ (.A1(_0548_),
    .A2(_0504_),
    .B(_0551_),
    .ZN(_0552_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5245_ (.I(_4336_),
    .Z(_0553_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _5246_ (.A1(_0544_),
    .A2(_0547_),
    .B1(_0552_),
    .B2(_0553_),
    .ZN(_0554_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5247_ (.I(_4315_),
    .Z(_0555_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _5248_ (.A1(_0549_),
    .A2(_0504_),
    .Z(_0556_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _5249_ (.A1(_0444_),
    .A2(_0453_),
    .B1(_0466_),
    .B2(_0442_),
    .ZN(_0557_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _5250_ (.A1(_0556_),
    .A2(_0557_),
    .Z(_0558_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5251_ (.A1(_0549_),
    .A2(_4421_),
    .ZN(_0559_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5252_ (.A1(_4488_),
    .A2(_0504_),
    .B(_0559_),
    .ZN(_0560_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5253_ (.I(_0560_),
    .Z(_0561_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5254_ (.I(_4338_),
    .Z(_0562_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _5255_ (.A1(_0555_),
    .A2(_0558_),
    .B1(_0561_),
    .B2(_0418_),
    .C(_0562_),
    .ZN(_0563_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5256_ (.A1(_0554_),
    .A2(_0563_),
    .ZN(_0564_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5257_ (.I(_0562_),
    .Z(_0565_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5258_ (.I(_0542_),
    .Z(_0566_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5259_ (.A1(\as2650.holding_reg[4] ),
    .A2(_0566_),
    .ZN(_0567_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _5260_ (.A1(_0565_),
    .A2(_0567_),
    .B(_0396_),
    .ZN(_0568_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_2 _5261_ (.A1(_0396_),
    .A2(_0543_),
    .B1(_0564_),
    .B2(_0568_),
    .ZN(_0569_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5262_ (.I(_0569_),
    .Z(_0570_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _5263_ (.I(_4502_),
    .Z(_0571_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _5264_ (.A1(_0477_),
    .A2(_0541_),
    .Z(_0572_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _5265_ (.A1(_4359_),
    .A2(_0503_),
    .Z(_0573_));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _5266_ (.A1(_0290_),
    .A2(_0481_),
    .A3(_0502_),
    .Z(_0574_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _5267_ (.A1(_0290_),
    .A2(_0481_),
    .B(_0502_),
    .ZN(_0575_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _5268_ (.A1(_0384_),
    .A2(_0574_),
    .A3(_0575_),
    .ZN(_0576_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_2 _5269_ (.A1(_0571_),
    .A2(_0572_),
    .B(_0573_),
    .C(_0576_),
    .ZN(_0577_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5270_ (.I(_0577_),
    .Z(_0578_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5271_ (.I(_0500_),
    .Z(_0579_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5272_ (.I(_0579_),
    .ZN(_0580_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _5273_ (.I0(\as2650.r123[1][5] ),
    .I1(\as2650.r123[0][5] ),
    .I2(\as2650.r123_2[1][5] ),
    .I3(\as2650.r123_2[0][5] ),
    .S0(_4196_),
    .S1(_0493_),
    .Z(_0581_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5274_ (.A1(_4521_),
    .A2(_0581_),
    .ZN(_0582_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _5275_ (.I0(\as2650.r123[2][5] ),
    .I1(\as2650.r123_2[2][5] ),
    .S(_0493_),
    .Z(_0583_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5276_ (.A1(_4298_),
    .A2(_0583_),
    .ZN(_0584_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5277_ (.I(\as2650.r0[5] ),
    .Z(_0585_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5278_ (.I(_0585_),
    .Z(_0586_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5279_ (.A1(_0586_),
    .A2(_4141_),
    .ZN(_0587_));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _5280_ (.A1(_0582_),
    .A2(_0584_),
    .A3(_0587_),
    .Z(_0588_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5281_ (.I(_0588_),
    .Z(_0589_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5282_ (.I(_0589_),
    .Z(_0590_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _5283_ (.I(_0590_),
    .Z(_0591_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5284_ (.I(_0591_),
    .Z(_0592_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5285_ (.I(_0592_),
    .Z(_0593_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5286_ (.I(net10),
    .Z(_0594_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5287_ (.I(_0594_),
    .Z(_0595_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5288_ (.I(_0595_),
    .Z(_0596_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5289_ (.I(_0596_),
    .Z(_0597_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5290_ (.I(_4396_),
    .Z(_0598_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5291_ (.A1(_4508_),
    .A2(_0480_),
    .ZN(_0599_));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _5292_ (.A1(_4182_),
    .A2(_4158_),
    .A3(_4177_),
    .Z(_0600_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5293_ (.A1(_4155_),
    .A2(_0600_),
    .ZN(_0601_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _5294_ (.A1(_0509_),
    .A2(_0463_),
    .B1(_0599_),
    .B2(_0601_),
    .ZN(_0602_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_2 _5295_ (.A1(_0503_),
    .A2(_0602_),
    .Z(_0603_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5296_ (.A1(_4397_),
    .A2(_0603_),
    .ZN(_0604_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _5297_ (.A1(_0597_),
    .A2(_0598_),
    .B(_0604_),
    .C(_4389_),
    .ZN(_0605_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _5298_ (.A1(_4378_),
    .A2(_0593_),
    .B(_0605_),
    .C(_4222_),
    .ZN(_0606_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _5299_ (.A1(_4364_),
    .A2(_0372_),
    .B(_0606_),
    .C(_4362_),
    .ZN(_0607_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _5300_ (.A1(_0580_),
    .A2(_4363_),
    .B(_4501_),
    .C(_0607_),
    .ZN(_0608_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _5301_ (.A1(_4501_),
    .A2(_0578_),
    .B(_0608_),
    .C(_0285_),
    .ZN(_0609_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _5302_ (.I(_4351_),
    .Z(_0610_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5303_ (.I(_4348_),
    .Z(_0611_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _5304_ (.A1(_0348_),
    .A2(_0574_),
    .A3(_0575_),
    .ZN(_0612_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_2 _5305_ (.A1(_0610_),
    .A2(_0503_),
    .B1(_0572_),
    .B2(_0611_),
    .C(_0612_),
    .ZN(_0613_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5306_ (.I(_0613_),
    .Z(_0614_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _5307_ (.A1(_4346_),
    .A2(_0614_),
    .B(_4412_),
    .ZN(_0615_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_2 _5308_ (.A1(_4276_),
    .A2(_0570_),
    .B1(_0609_),
    .B2(_0615_),
    .ZN(_0616_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5309_ (.I(_0580_),
    .Z(_0617_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5310_ (.I(_4426_),
    .Z(_0618_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5311_ (.I(_0618_),
    .Z(_0619_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5312_ (.I(_0619_),
    .Z(_0620_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5313_ (.I(_0620_),
    .Z(_0621_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5314_ (.I(_4452_),
    .Z(_0622_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5315_ (.A1(\as2650.stack[3][12] ),
    .A2(_0622_),
    .B(_4454_),
    .ZN(_0623_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5316_ (.I(_4460_),
    .Z(_0624_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5317_ (.A1(\as2650.stack[2][12] ),
    .A2(_0624_),
    .ZN(_0625_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5318_ (.I(_0324_),
    .Z(_0626_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _5319_ (.A1(\as2650.stack[0][12] ),
    .A2(_4482_),
    .B1(_0626_),
    .B2(\as2650.stack[1][12] ),
    .ZN(_0627_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _5320_ (.A1(_0623_),
    .A2(_0625_),
    .A3(_0627_),
    .ZN(_0628_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _5321_ (.A1(\as2650.stack[4][12] ),
    .A2(_4482_),
    .B1(_0626_),
    .B2(\as2650.stack[5][12] ),
    .ZN(_0629_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _5322_ (.A1(\as2650.stack[7][12] ),
    .A2(_4479_),
    .B1(_4461_),
    .B2(\as2650.stack[6][12] ),
    .ZN(_0630_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _5323_ (.A1(_4477_),
    .A2(_0629_),
    .A3(_0630_),
    .ZN(_0631_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5324_ (.A1(_0628_),
    .A2(_0631_),
    .ZN(_0632_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _5325_ (.A1(_0617_),
    .A2(_0621_),
    .B1(_4446_),
    .B2(_0632_),
    .C(_0438_),
    .ZN(_0633_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _5326_ (.A1(_4500_),
    .A2(_0616_),
    .B(_0633_),
    .C(_0538_),
    .ZN(_0634_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _5327_ (.A1(_0540_),
    .A2(_4499_),
    .B(_0634_),
    .ZN(_0004_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5328_ (.I(\as2650.r123[0][5] ),
    .ZN(_0635_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5329_ (.I(_0395_),
    .Z(_0636_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5330_ (.I(\as2650.holding_reg[5] ),
    .Z(_0637_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _5331_ (.A1(_0582_),
    .A2(_0584_),
    .A3(_0587_),
    .ZN(_0638_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5332_ (.I(_0638_),
    .Z(_0639_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _5333_ (.A1(_0637_),
    .A2(_0639_),
    .Z(_0640_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5334_ (.I(_0640_),
    .Z(_0641_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _5335_ (.A1(\as2650.holding_reg[5] ),
    .A2(_0591_),
    .Z(_0642_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5336_ (.I(_0567_),
    .ZN(_0643_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _5337_ (.A1(_0543_),
    .A2(_0546_),
    .B(_0643_),
    .ZN(_0644_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _5338_ (.A1(_0642_),
    .A2(_0644_),
    .Z(_0645_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5339_ (.A1(_0544_),
    .A2(_0645_),
    .ZN(_0646_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _5340_ (.A1(_0556_),
    .A2(_0557_),
    .B1(_0560_),
    .B2(_0567_),
    .ZN(_0647_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5341_ (.A1(_0641_),
    .A2(_0647_),
    .ZN(_0648_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _5342_ (.A1(_0640_),
    .A2(_0647_),
    .Z(_0649_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _5343_ (.A1(_0555_),
    .A2(_0648_),
    .A3(_0649_),
    .ZN(_0650_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5344_ (.I(_0418_),
    .Z(_0651_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5345_ (.A1(\as2650.holding_reg[5] ),
    .A2(_4191_),
    .ZN(_0652_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _5346_ (.A1(_4421_),
    .A2(_0591_),
    .B(_0652_),
    .ZN(_0653_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5347_ (.I(_0414_),
    .Z(_0654_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5348_ (.A1(_0637_),
    .A2(_0548_),
    .ZN(_0655_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5349_ (.A1(_0654_),
    .A2(_0592_),
    .B(_0655_),
    .ZN(_0656_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _5350_ (.A1(_0651_),
    .A2(_0653_),
    .B1(_0656_),
    .B2(_0553_),
    .C(_0562_),
    .ZN(_0657_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _5351_ (.A1(_0646_),
    .A2(_0650_),
    .A3(_0657_),
    .ZN(_0658_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5352_ (.A1(_0637_),
    .A2(_0638_),
    .ZN(_0659_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _5353_ (.A1(_0565_),
    .A2(_0659_),
    .B(_0396_),
    .ZN(_0660_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _5354_ (.A1(_0636_),
    .A2(_0641_),
    .B1(_0658_),
    .B2(_0660_),
    .ZN(_0661_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5355_ (.I(_0661_),
    .Z(_0662_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _5356_ (.A1(_0589_),
    .A2(_0574_),
    .Z(_0663_));
 gf180mcu_fd_sc_mcu7t5v0__and4_1 _5357_ (.A1(_0349_),
    .A2(_4505_),
    .A3(_0369_),
    .A4(_0541_),
    .Z(_0664_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _5358_ (.A1(_0589_),
    .A2(_0664_),
    .Z(_0665_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _5359_ (.A1(_0611_),
    .A2(_0665_),
    .Z(_0666_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_2 _5360_ (.A1(_0610_),
    .A2(_0590_),
    .B1(_0663_),
    .B2(_4350_),
    .C(_0666_),
    .ZN(_0667_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5361_ (.I(_0667_),
    .Z(_0668_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5362_ (.I(_0586_),
    .Z(_0669_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5363_ (.I(_0669_),
    .Z(_0670_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5364_ (.I(\as2650.r0[6] ),
    .Z(_0671_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5365_ (.I(_0671_),
    .Z(_0672_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5366_ (.A1(_0672_),
    .A2(_4142_),
    .ZN(_0673_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _5367_ (.I0(\as2650.r123[2][6] ),
    .I1(\as2650.r123_2[2][6] ),
    .S(_0493_),
    .Z(_0674_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5368_ (.A1(_4369_),
    .A2(_0674_),
    .ZN(_0675_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _5369_ (.I0(\as2650.r123[1][6] ),
    .I1(\as2650.r123[0][6] ),
    .I2(\as2650.r123_2[1][6] ),
    .I3(\as2650.r123_2[0][6] ),
    .S0(_4196_),
    .S1(_4148_),
    .Z(_0676_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5370_ (.A1(_4300_),
    .A2(_0676_),
    .ZN(_0677_));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _5371_ (.A1(_0673_),
    .A2(_0675_),
    .A3(_0677_),
    .Z(_0678_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _5372_ (.I(_0678_),
    .Z(_0679_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5373_ (.I(_0679_),
    .Z(_0680_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5374_ (.I(_0680_),
    .Z(_0681_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5375_ (.I(net1),
    .Z(_0682_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5376_ (.I(_0682_),
    .Z(_0683_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5377_ (.I(_0683_),
    .Z(_0684_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5378_ (.I(_0684_),
    .Z(_0685_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_2 _5379_ (.A1(_0354_),
    .A2(_4506_),
    .A3(_0370_),
    .A4(_0542_),
    .ZN(_0686_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _5380_ (.A1(_4182_),
    .A2(_4193_),
    .ZN(_0687_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5381_ (.A1(_4155_),
    .A2(_0687_),
    .ZN(_0688_));
 gf180mcu_fd_sc_mcu7t5v0__oai32_1 _5382_ (.A1(_0601_),
    .A2(_0599_),
    .A3(_0542_),
    .B1(_0686_),
    .B2(_0688_),
    .ZN(_0689_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_2 _5383_ (.A1(_0590_),
    .A2(_0689_),
    .Z(_0690_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5384_ (.A1(_0598_),
    .A2(_0690_),
    .ZN(_0691_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _5385_ (.A1(_0685_),
    .A2(_4532_),
    .B(_0691_),
    .C(_4378_),
    .ZN(_0692_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _5386_ (.A1(_4515_),
    .A2(_0681_),
    .B(_0692_),
    .C(_4538_),
    .ZN(_0693_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5387_ (.I(_0505_),
    .Z(_0694_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _5388_ (.A1(_0517_),
    .A2(_0694_),
    .B(_4546_),
    .ZN(_0695_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _5389_ (.A1(_0670_),
    .A2(_4547_),
    .B1(_0693_),
    .B2(_0695_),
    .ZN(_0696_));
 gf180mcu_fd_sc_mcu7t5v0__aoi222_2 _5390_ (.A1(_0571_),
    .A2(_0665_),
    .B1(_0663_),
    .B2(_4358_),
    .C1(_0487_),
    .C2(_0591_),
    .ZN(_0697_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5391_ (.I(_0697_),
    .Z(_0698_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5392_ (.A1(_0486_),
    .A2(_0698_),
    .ZN(_0699_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5393_ (.I(_0284_),
    .Z(_0700_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _5394_ (.A1(_4354_),
    .A2(_0696_),
    .B(_0699_),
    .C(_0700_),
    .ZN(_0701_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _5395_ (.A1(_0285_),
    .A2(_0668_),
    .B(_0701_),
    .C(_0295_),
    .ZN(_0702_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5396_ (.A1(_0296_),
    .A2(_0662_),
    .B(_0702_),
    .ZN(_0703_));
 gf180mcu_fd_sc_mcu7t5v0__aoi222_2 _5397_ (.A1(\as2650.stack[7][13] ),
    .A2(_0326_),
    .B1(_4466_),
    .B2(\as2650.stack[4][13] ),
    .C1(\as2650.stack[5][13] ),
    .C2(_4470_),
    .ZN(_0704_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _5398_ (.A1(\as2650.stack[6][13] ),
    .A2(_4461_),
    .B(_0329_),
    .ZN(_0705_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _5399_ (.A1(\as2650.stack[0][13] ),
    .A2(_4481_),
    .B1(_0324_),
    .B2(\as2650.stack[1][13] ),
    .ZN(_0706_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5400_ (.I(_0706_),
    .ZN(_0707_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_2 _5401_ (.A1(\as2650.stack[3][13] ),
    .A2(_4479_),
    .B1(_0427_),
    .B2(\as2650.stack[2][13] ),
    .C(_0707_),
    .ZN(_0708_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_2 _5402_ (.A1(_0704_),
    .A2(_0705_),
    .B1(_0708_),
    .B2(_0526_),
    .ZN(_0709_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5403_ (.A1(_4485_),
    .A2(_0709_),
    .ZN(_0710_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5404_ (.I(_0670_),
    .Z(_0711_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5405_ (.A1(_0711_),
    .A2(_0343_),
    .ZN(_0712_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _5406_ (.A1(_0438_),
    .A2(_0710_),
    .A3(_0712_),
    .ZN(_0713_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _5407_ (.A1(_4274_),
    .A2(_0703_),
    .B(_0713_),
    .C(_0538_),
    .ZN(_0714_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _5408_ (.A1(_0635_),
    .A2(_4440_),
    .B(_0714_),
    .ZN(_0005_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5409_ (.I(\as2650.r123[0][6] ),
    .ZN(_0715_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _5410_ (.A1(_0673_),
    .A2(_0675_),
    .A3(_0677_),
    .ZN(_0716_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5411_ (.I(_0716_),
    .Z(_0717_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5412_ (.I(_0717_),
    .Z(_0718_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _5413_ (.A1(\as2650.holding_reg[6] ),
    .A2(_0718_),
    .Z(_0719_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5414_ (.I(_0719_),
    .Z(_0720_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5415_ (.I(_0719_),
    .ZN(_0721_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5416_ (.A1(_0659_),
    .A2(_0653_),
    .ZN(_0722_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5417_ (.A1(_0640_),
    .A2(_0647_),
    .B(_0722_),
    .ZN(_0723_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5418_ (.A1(_0721_),
    .A2(_0723_),
    .ZN(_0724_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _5419_ (.A1(_0649_),
    .A2(_0720_),
    .A3(_0722_),
    .ZN(_0725_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _5420_ (.A1(_0555_),
    .A2(_0724_),
    .A3(_0725_),
    .ZN(_0726_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5421_ (.A1(_0642_),
    .A2(_0644_),
    .B(_0659_),
    .ZN(_0727_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _5422_ (.A1(_0719_),
    .A2(_0727_),
    .B(_0411_),
    .ZN(_0728_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5423_ (.A1(_0720_),
    .A2(_0727_),
    .B(_0728_),
    .ZN(_0729_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5424_ (.I(\as2650.holding_reg[6] ),
    .Z(_0730_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5425_ (.A1(_0730_),
    .A2(_0469_),
    .ZN(_0731_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _5426_ (.A1(_4427_),
    .A2(_0679_),
    .B(_0731_),
    .ZN(_0732_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5427_ (.A1(_0730_),
    .A2(_0548_),
    .ZN(_0733_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5428_ (.A1(_0654_),
    .A2(_0680_),
    .B(_0733_),
    .ZN(_0734_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _5429_ (.A1(_0651_),
    .A2(_0732_),
    .B1(_0734_),
    .B2(_0553_),
    .C(_0562_),
    .ZN(_0735_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _5430_ (.A1(_0726_),
    .A2(_0729_),
    .A3(_0735_),
    .ZN(_0736_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5431_ (.A1(_0730_),
    .A2(_0718_),
    .ZN(_0737_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _5432_ (.A1(_0565_),
    .A2(_0737_),
    .B(_0636_),
    .ZN(_0738_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _5433_ (.A1(_0636_),
    .A2(_0720_),
    .B1(_0736_),
    .B2(_0738_),
    .ZN(_0739_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5434_ (.I(_0739_),
    .Z(_0740_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _5435_ (.A1(_0638_),
    .A2(_0664_),
    .A3(_0716_),
    .ZN(_0741_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5436_ (.A1(_0590_),
    .A2(_0686_),
    .B(_0678_),
    .ZN(_0742_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5437_ (.A1(_0741_),
    .A2(_0742_),
    .ZN(_0743_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5438_ (.A1(_0502_),
    .A2(_0588_),
    .ZN(_0744_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5439_ (.A1(_0599_),
    .A2(_0744_),
    .ZN(_0745_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _5440_ (.A1(_0745_),
    .A2(_0716_),
    .Z(_0746_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5441_ (.A1(_0348_),
    .A2(_0746_),
    .ZN(_0747_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_2 _5442_ (.A1(_0610_),
    .A2(_0678_),
    .B1(_0743_),
    .B2(_0611_),
    .C(_0747_),
    .ZN(_0748_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5443_ (.I(_0748_),
    .Z(_0749_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5444_ (.I(_0672_),
    .Z(_0750_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5445_ (.I(_0750_),
    .Z(_0751_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5446_ (.I(_0751_),
    .Z(_0752_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5447_ (.I(_4376_),
    .Z(_0753_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5448_ (.I(_0753_),
    .Z(_0754_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5449_ (.I(net2),
    .Z(_0755_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5450_ (.I(_0755_),
    .Z(_0756_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5451_ (.I(_0756_),
    .Z(_0757_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5452_ (.I(_0757_),
    .Z(_0758_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5453_ (.I(_0758_),
    .Z(_0759_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _5454_ (.A1(_4533_),
    .A2(_0589_),
    .A3(_0574_),
    .ZN(_0760_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _5455_ (.A1(_4218_),
    .A2(_0638_),
    .A3(_0664_),
    .ZN(_0761_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5456_ (.A1(_0760_),
    .A2(_0761_),
    .ZN(_0762_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _5457_ (.A1(_0679_),
    .A2(_0762_),
    .Z(_0763_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5458_ (.A1(_0598_),
    .A2(_0763_),
    .ZN(_0764_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _5459_ (.A1(_0759_),
    .A2(_4532_),
    .B(_0764_),
    .C(_4231_),
    .ZN(_0765_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _5460_ (.A1(_4515_),
    .A2(_0754_),
    .B(_0765_),
    .C(_4538_),
    .ZN(_0766_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _5461_ (.A1(_0517_),
    .A2(_0593_),
    .B(_4546_),
    .ZN(_0767_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _5462_ (.A1(_0752_),
    .A2(_4547_),
    .B1(_0766_),
    .B2(_0767_),
    .ZN(_0768_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5463_ (.A1(_0384_),
    .A2(_0746_),
    .ZN(_0769_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_2 _5464_ (.A1(_0487_),
    .A2(_0679_),
    .B1(_0743_),
    .B2(_0571_),
    .C(_0769_),
    .ZN(_0770_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5465_ (.I(_0770_),
    .Z(_0771_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5466_ (.A1(_0486_),
    .A2(_0771_),
    .ZN(_0772_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _5467_ (.A1(_4354_),
    .A2(_0768_),
    .B(_0772_),
    .C(_0700_),
    .ZN(_0773_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _5468_ (.A1(_0285_),
    .A2(_0749_),
    .B(_0773_),
    .C(_0295_),
    .ZN(_0774_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _5469_ (.A1(_0296_),
    .A2(_0740_),
    .B(_0774_),
    .ZN(_0775_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _5470_ (.A1(\as2650.stack[7][14] ),
    .A2(_0326_),
    .B1(_0527_),
    .B2(\as2650.stack[6][14] ),
    .ZN(_0776_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_2 _5471_ (.A1(\as2650.stack[4][14] ),
    .A2(_4481_),
    .B1(_0430_),
    .B2(\as2650.stack[5][14] ),
    .C(_0329_),
    .ZN(_0777_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _5472_ (.A1(\as2650.stack[0][14] ),
    .A2(_4465_),
    .B1(_4469_),
    .B2(\as2650.stack[1][14] ),
    .ZN(_0778_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5473_ (.I(_0778_),
    .ZN(_0779_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_2 _5474_ (.A1(\as2650.stack[3][14] ),
    .A2(_4478_),
    .B1(_0527_),
    .B2(\as2650.stack[2][14] ),
    .C(_0779_),
    .ZN(_0780_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_2 _5475_ (.A1(_0776_),
    .A2(_0777_),
    .B1(_0780_),
    .B2(_0526_),
    .ZN(_0781_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5476_ (.A1(_4445_),
    .A2(_0781_),
    .ZN(_0782_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5477_ (.A1(_0752_),
    .A2(_0343_),
    .ZN(_0783_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _5478_ (.A1(_0438_),
    .A2(_0782_),
    .A3(_0783_),
    .ZN(_0784_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _5479_ (.A1(_4274_),
    .A2(_0775_),
    .B(_0784_),
    .C(_0538_),
    .ZN(_0785_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _5480_ (.A1(_0715_),
    .A2(_4440_),
    .B(_0785_),
    .ZN(_0006_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5481_ (.I(\as2650.r123[0][7] ),
    .ZN(_0786_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5482_ (.I(_4494_),
    .ZN(_0787_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5483_ (.I(_4367_),
    .Z(_0788_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5484_ (.I(_0788_),
    .Z(_0789_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5485_ (.I(_0789_),
    .Z(_0790_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5486_ (.I(_0790_),
    .Z(_0791_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _5487_ (.A1(_0791_),
    .A2(_0620_),
    .Z(_0792_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _5488_ (.A1(_0787_),
    .A2(_0792_),
    .B(_4498_),
    .ZN(_0793_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _5489_ (.A1(\as2650.holding_reg[7] ),
    .A2(_4376_),
    .Z(_0794_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5490_ (.I(_0794_),
    .Z(_0795_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _5491_ (.A1(_0721_),
    .A2(_0723_),
    .Z(_0796_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5492_ (.A1(_0737_),
    .A2(_0732_),
    .ZN(_0797_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5493_ (.I(_0797_),
    .ZN(_0798_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _5494_ (.A1(_4368_),
    .A2(_4371_),
    .A3(_4373_),
    .ZN(_0799_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _5495_ (.A1(\as2650.holding_reg[7] ),
    .A2(_0799_),
    .Z(_0800_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _5496_ (.I(_0800_),
    .Z(_0801_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5497_ (.A1(_0796_),
    .A2(_0798_),
    .B(_0801_),
    .ZN(_0802_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _5498_ (.A1(_0724_),
    .A2(_0794_),
    .A3(_0797_),
    .ZN(_0803_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _5499_ (.A1(_0802_),
    .A2(_0803_),
    .B(_0448_),
    .ZN(_0804_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5500_ (.I(_0737_),
    .ZN(_0805_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _5501_ (.A1(_0719_),
    .A2(_0727_),
    .B(_0805_),
    .ZN(_0806_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _5502_ (.A1(_0794_),
    .A2(_0806_),
    .Z(_0807_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _5503_ (.A1(_0544_),
    .A2(_0807_),
    .Z(_0808_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5504_ (.A1(\as2650.holding_reg[7] ),
    .A2(_0550_),
    .ZN(_0809_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5505_ (.A1(_0550_),
    .A2(_4376_),
    .B(_0809_),
    .ZN(_0810_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5506_ (.A1(_4336_),
    .A2(_0810_),
    .ZN(_0811_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5507_ (.A1(_0313_),
    .A2(_0811_),
    .ZN(_0812_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5508_ (.I(\as2650.holding_reg[7] ),
    .Z(_0813_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5509_ (.I(_0447_),
    .Z(_0814_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5510_ (.A1(_0813_),
    .A2(_0799_),
    .B(_0814_),
    .ZN(_0815_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5511_ (.A1(_0651_),
    .A2(_0815_),
    .ZN(_0816_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_1 _5512_ (.A1(_0804_),
    .A2(_0808_),
    .A3(_0812_),
    .B(_0816_),
    .ZN(_0817_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5513_ (.I(_0799_),
    .Z(_0818_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _5514_ (.A1(_0813_),
    .A2(_0565_),
    .A3(_0818_),
    .ZN(_0819_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _5515_ (.A1(_0473_),
    .A2(_0819_),
    .Z(_0820_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_2 _5516_ (.A1(_0636_),
    .A2(_0795_),
    .B1(_0817_),
    .B2(_0820_),
    .ZN(_0821_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _5517_ (.A1(_0799_),
    .A2(_0741_),
    .Z(_0822_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5518_ (.A1(_0611_),
    .A2(_0822_),
    .ZN(_0823_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_2 _5519_ (.A1(_0599_),
    .A2(_0744_),
    .A3(_0717_),
    .ZN(_0824_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _5520_ (.A1(_4374_),
    .A2(_0824_),
    .Z(_0825_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _5521_ (.A1(_4375_),
    .A2(_0610_),
    .B1(_0825_),
    .B2(_4350_),
    .ZN(_0826_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5522_ (.A1(_0823_),
    .A2(_0826_),
    .ZN(_0827_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5523_ (.I(_0827_),
    .Z(_0828_));
 gf180mcu_fd_sc_mcu7t5v0__aoi222_2 _5524_ (.A1(_4375_),
    .A2(_0487_),
    .B1(_0822_),
    .B2(_0571_),
    .C1(_0825_),
    .C2(_4358_),
    .ZN(_0829_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5525_ (.I(_0829_),
    .Z(_0830_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5526_ (.A1(_4408_),
    .A2(_0830_),
    .B(_0700_),
    .ZN(_0831_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _5527_ (.I0(_0760_),
    .I1(_0761_),
    .S(_0717_),
    .Z(_0832_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _5528_ (.A1(_4375_),
    .A2(_0832_),
    .Z(_0833_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5529_ (.I(_0833_),
    .Z(_0834_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5530_ (.I(net3),
    .ZN(_0835_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5531_ (.I(_0835_),
    .Z(_0836_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _5532_ (.I(_0836_),
    .Z(_0837_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5533_ (.A1(_0837_),
    .A2(_0598_),
    .B(_4231_),
    .ZN(_0838_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _5534_ (.A1(_4532_),
    .A2(_0834_),
    .B(_0838_),
    .ZN(_0839_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5535_ (.A1(_4320_),
    .A2(_4334_),
    .B(_4321_),
    .ZN(_0840_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5536_ (.A1(_4515_),
    .A2(_0840_),
    .ZN(_0841_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5537_ (.A1(_0839_),
    .A2(_0841_),
    .B(_4364_),
    .ZN(_0842_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _5538_ (.A1(_0517_),
    .A2(_0681_),
    .B(_4546_),
    .ZN(_0843_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _5539_ (.A1(_0790_),
    .A2(_4547_),
    .B1(_0842_),
    .B2(_0843_),
    .C(_0486_),
    .ZN(_0844_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_1 _5540_ (.A1(_0700_),
    .A2(_0828_),
    .B1(_0831_),
    .B2(_0844_),
    .C(_0295_),
    .ZN(_0845_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5541_ (.A1(_0296_),
    .A2(_0821_),
    .B(_0845_),
    .ZN(_0846_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _5542_ (.A1(_4275_),
    .A2(_0846_),
    .Z(_0847_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _5543_ (.A1(_0786_),
    .A2(_4440_),
    .B1(_0793_),
    .B2(_0847_),
    .ZN(_0007_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5544_ (.I(_4295_),
    .Z(_0848_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5545_ (.I(_4448_),
    .Z(_0849_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5546_ (.I(_0849_),
    .Z(_0850_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5547_ (.I(_0850_),
    .Z(_0851_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _5548_ (.I(_4204_),
    .Z(_0852_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5549_ (.I(_4487_),
    .Z(_0853_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _5550_ (.A1(_4488_),
    .A2(_4429_),
    .A3(_4424_),
    .ZN(_0854_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _5551_ (.A1(_0853_),
    .A2(_0854_),
    .Z(_0855_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5552_ (.A1(_0852_),
    .A2(_0855_),
    .ZN(_0856_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5553_ (.I(_0856_),
    .Z(_0857_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5554_ (.I(_0857_),
    .Z(_0858_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _5555_ (.A1(_0851_),
    .A2(_0626_),
    .A3(_0858_),
    .ZN(_0859_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _5556_ (.I(_0859_),
    .Z(_0860_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5557_ (.I(_0860_),
    .Z(_0861_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5558_ (.I(\as2650.pc[0] ),
    .Z(_0862_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5559_ (.I(_0862_),
    .ZN(_0863_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5560_ (.I(_0863_),
    .Z(_0864_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5561_ (.I(_0864_),
    .Z(_0865_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5562_ (.I(_0850_),
    .Z(_0866_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5563_ (.I(_4214_),
    .Z(_0867_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5564_ (.I(_4215_),
    .Z(_0868_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _5565_ (.A1(_4224_),
    .A2(_4369_),
    .A3(_4313_),
    .ZN(_0869_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5566_ (.A1(_4255_),
    .A2(_0869_),
    .ZN(_0870_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5567_ (.I(_0870_),
    .Z(_0871_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5568_ (.A1(_0868_),
    .A2(_0871_),
    .ZN(_0872_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5569_ (.A1(_0867_),
    .A2(_0872_),
    .ZN(_0873_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5570_ (.I(_4184_),
    .Z(_0874_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5571_ (.A1(_0874_),
    .A2(_4193_),
    .ZN(_0875_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5572_ (.I(_4180_),
    .Z(_0876_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5573_ (.I(_0876_),
    .Z(_0877_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5574_ (.A1(_4207_),
    .A2(_4175_),
    .ZN(_0878_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5575_ (.I(_0878_),
    .Z(_0879_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5576_ (.A1(_0877_),
    .A2(_0879_),
    .ZN(_0880_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5577_ (.I(\as2650.addr_buff[7] ),
    .Z(_0881_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5578_ (.I(_4254_),
    .Z(_0882_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5579_ (.I(_4208_),
    .Z(_0883_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5580_ (.I(\as2650.cycle[1] ),
    .Z(_0884_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5581_ (.I(_4238_),
    .ZN(_0885_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _5582_ (.I(_4239_),
    .Z(_0886_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _5583_ (.A1(_4234_),
    .A2(_0885_),
    .A3(_0886_),
    .ZN(_0887_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_2 _5584_ (.A1(_4251_),
    .A2(_4164_),
    .A3(_0884_),
    .A4(_0887_),
    .ZN(_0888_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5585_ (.A1(_0883_),
    .A2(_0888_),
    .ZN(_0889_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5586_ (.A1(_0881_),
    .A2(_0882_),
    .B(_0889_),
    .ZN(_0890_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5587_ (.A1(_0877_),
    .A2(_0870_),
    .ZN(_0891_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _5588_ (.A1(_0836_),
    .A2(_0880_),
    .B1(_0890_),
    .B2(_0891_),
    .ZN(_0892_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _5589_ (.I(_4251_),
    .Z(_0893_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _5590_ (.A1(_0893_),
    .A2(_4164_),
    .A3(_4172_),
    .ZN(_0894_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _5591_ (.A1(_0884_),
    .A2(_4208_),
    .A3(_0894_),
    .ZN(_0895_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5592_ (.I(_0895_),
    .Z(_0896_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5593_ (.A1(_0447_),
    .A2(_0896_),
    .ZN(_0897_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5594_ (.I(_0891_),
    .Z(_0898_));
 gf180mcu_fd_sc_mcu7t5v0__oai32_1 _5595_ (.A1(_0873_),
    .A2(_0875_),
    .A3(_0892_),
    .B1(_0897_),
    .B2(_0898_),
    .ZN(_0899_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _5596_ (.A1(_4152_),
    .A2(_0899_),
    .Z(_0900_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5597_ (.I(_0900_),
    .Z(_0901_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _5598_ (.A1(_0866_),
    .A2(_4466_),
    .A3(_0901_),
    .ZN(_0902_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5599_ (.I(_0902_),
    .Z(_0903_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5600_ (.I(_0902_),
    .Z(_0904_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5601_ (.A1(\as2650.stack[5][0] ),
    .A2(_0904_),
    .ZN(_0905_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5602_ (.A1(_0865_),
    .A2(_0903_),
    .B(_0905_),
    .ZN(_0906_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5603_ (.A1(_0861_),
    .A2(_0906_),
    .ZN(_0907_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5604_ (.A1(_0848_),
    .A2(_0861_),
    .B(_0907_),
    .ZN(_0008_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5605_ (.I(_0337_),
    .Z(_0908_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5606_ (.I(\as2650.pc[1] ),
    .Z(_0909_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5607_ (.I(_0909_),
    .Z(_0910_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5608_ (.I(_0910_),
    .Z(_0911_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5609_ (.I(_0911_),
    .Z(_0912_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5610_ (.I(_0902_),
    .Z(_0913_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _5611_ (.I0(_0912_),
    .I1(\as2650.stack[5][1] ),
    .S(_0913_),
    .Z(_0914_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _5612_ (.I(_0859_),
    .Z(_0915_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _5613_ (.I0(_0908_),
    .I1(_0914_),
    .S(_0915_),
    .Z(_0916_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5614_ (.I(_0916_),
    .Z(_0009_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5615_ (.I(_0361_),
    .Z(_0917_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5616_ (.I(_0917_),
    .Z(_0918_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5617_ (.I(\as2650.pc[2] ),
    .Z(_0919_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5618_ (.I(_0919_),
    .Z(_0920_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5619_ (.I(_0920_),
    .Z(_0921_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _5620_ (.I0(_0921_),
    .I1(\as2650.stack[5][2] ),
    .S(_0913_),
    .Z(_0922_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _5621_ (.I0(_0918_),
    .I1(_0922_),
    .S(_0915_),
    .Z(_0923_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5622_ (.I(_0923_),
    .Z(_0010_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5623_ (.I(_0535_),
    .Z(_0924_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5624_ (.I(_0924_),
    .Z(_0925_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5625_ (.I(\as2650.pc[3] ),
    .ZN(_0926_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5626_ (.I(_0926_),
    .Z(_0927_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5627_ (.I(_0927_),
    .Z(_0928_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5628_ (.A1(\as2650.stack[5][3] ),
    .A2(_0904_),
    .ZN(_0929_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5629_ (.A1(_0928_),
    .A2(_0903_),
    .B(_0929_),
    .ZN(_0930_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _5630_ (.I0(_0925_),
    .I1(_0930_),
    .S(_0860_),
    .Z(_0931_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5631_ (.I(_0931_),
    .Z(_0011_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5632_ (.I(_0617_),
    .Z(_0932_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _5633_ (.I(\as2650.pc[4] ),
    .ZN(_0933_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5634_ (.A1(\as2650.stack[5][4] ),
    .A2(_0913_),
    .ZN(_0934_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5635_ (.A1(_0933_),
    .A2(_0903_),
    .B(_0934_),
    .ZN(_0935_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5636_ (.A1(_0915_),
    .A2(_0935_),
    .ZN(_0936_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5637_ (.A1(_0932_),
    .A2(_0861_),
    .B(_0936_),
    .ZN(_0012_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5638_ (.I(_0711_),
    .ZN(_0937_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5639_ (.I(_0937_),
    .Z(_0938_));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _5640_ (.I(\as2650.pc[5] ),
    .ZN(_0939_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5641_ (.I(_0939_),
    .Z(_0940_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5642_ (.A1(\as2650.stack[5][5] ),
    .A2(_0913_),
    .ZN(_0941_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5643_ (.A1(_0940_),
    .A2(_0904_),
    .B(_0941_),
    .ZN(_0942_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5644_ (.A1(_0915_),
    .A2(_0942_),
    .ZN(_0943_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5645_ (.A1(_0938_),
    .A2(_0861_),
    .B(_0943_),
    .ZN(_0013_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5646_ (.I(_0752_),
    .Z(_0944_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5647_ (.I(\as2650.pc[6] ),
    .Z(_0945_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5648_ (.I(_0945_),
    .Z(_0946_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5649_ (.I(_0946_),
    .Z(_0947_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5650_ (.I(_0947_),
    .Z(_0948_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _5651_ (.I0(_0948_),
    .I1(\as2650.stack[5][6] ),
    .S(_0902_),
    .Z(_0949_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _5652_ (.I0(_0944_),
    .I1(_0949_),
    .S(_0860_),
    .Z(_0950_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5653_ (.I(_0950_),
    .Z(_0014_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5654_ (.I(_0791_),
    .Z(_0951_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5655_ (.I(\as2650.pc[7] ),
    .ZN(_0952_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5656_ (.I(_0952_),
    .Z(_0953_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5657_ (.A1(\as2650.stack[5][7] ),
    .A2(_0904_),
    .ZN(_0954_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5658_ (.A1(_0953_),
    .A2(_0903_),
    .B(_0954_),
    .ZN(_0955_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _5659_ (.I0(_0951_),
    .I1(_0955_),
    .S(_0860_),
    .Z(_0956_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5660_ (.I(_0956_),
    .Z(_0015_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5661_ (.I(_0850_),
    .Z(_0957_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5662_ (.A1(_0957_),
    .A2(_0430_),
    .ZN(_0958_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5663_ (.A1(_0856_),
    .A2(_0900_),
    .ZN(_0959_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5664_ (.I(_0959_),
    .Z(_0960_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5665_ (.A1(_0958_),
    .A2(_0960_),
    .ZN(_0961_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5666_ (.I(_0961_),
    .Z(_0962_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5667_ (.I(_0962_),
    .Z(_0963_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5668_ (.I(\as2650.pc[8] ),
    .Z(_0964_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5669_ (.I(_0964_),
    .Z(_0965_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5670_ (.I(_0965_),
    .Z(_0966_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5671_ (.I(_0857_),
    .Z(_0967_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5672_ (.I(_0967_),
    .Z(_0968_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5673_ (.I(_4152_),
    .Z(_0969_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5674_ (.A1(_4487_),
    .A2(_0854_),
    .ZN(_0970_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5675_ (.I(_0970_),
    .Z(_0971_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _5676_ (.A1(_0294_),
    .A2(_0969_),
    .A3(_0971_),
    .ZN(_0972_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _5677_ (.I(_0972_),
    .Z(_0973_));
 gf180mcu_fd_sc_mcu7t5v0__or3_1 _5678_ (.A1(\as2650.r123[0][0] ),
    .A2(_4153_),
    .A3(_0855_),
    .Z(_0974_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_1 _5679_ (.A1(_0966_),
    .A2(_0968_),
    .B1(_0973_),
    .B2(\as2650.r123_2[0][0] ),
    .C(_0974_),
    .ZN(_0975_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5680_ (.I(_0975_),
    .Z(_0976_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5681_ (.I(_0962_),
    .Z(_0977_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5682_ (.A1(\as2650.stack[6][8] ),
    .A2(_0977_),
    .ZN(_0978_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _5683_ (.A1(_0963_),
    .A2(_0976_),
    .B(_0978_),
    .ZN(_0016_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5684_ (.I(\as2650.pc[9] ),
    .Z(_0979_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _5685_ (.I(_0967_),
    .Z(_0980_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5686_ (.I(_4415_),
    .Z(_0981_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5687_ (.I(_0971_),
    .Z(_0982_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _5688_ (.A1(_4497_),
    .A2(_0981_),
    .A3(_0982_),
    .ZN(_0983_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_2 _5689_ (.A1(_0979_),
    .A2(_0980_),
    .B1(_0973_),
    .B2(\as2650.r123_2[0][1] ),
    .C(_0983_),
    .ZN(_0984_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5690_ (.I(_0984_),
    .Z(_0985_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5691_ (.I(_0961_),
    .Z(_0986_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5692_ (.A1(\as2650.stack[6][9] ),
    .A2(_0986_),
    .ZN(_0987_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _5693_ (.A1(_0963_),
    .A2(_0985_),
    .B(_0987_),
    .ZN(_0017_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5694_ (.I(\as2650.pc[10] ),
    .Z(_0988_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5695_ (.I(_0988_),
    .Z(_0989_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5696_ (.I(_0989_),
    .Z(_0990_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _5697_ (.A1(_0347_),
    .A2(_0981_),
    .A3(_0982_),
    .ZN(_0991_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_2 _5698_ (.A1(_0990_),
    .A2(_0980_),
    .B1(_0973_),
    .B2(\as2650.r123_2[0][2] ),
    .C(_0991_),
    .ZN(_0992_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5699_ (.I(_0992_),
    .Z(_0993_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5700_ (.A1(\as2650.stack[6][10] ),
    .A2(_0986_),
    .ZN(_0994_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _5701_ (.A1(_0963_),
    .A2(_0993_),
    .B(_0994_),
    .ZN(_0018_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5702_ (.I(\as2650.pc[11] ),
    .Z(_0995_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5703_ (.I(_0995_),
    .Z(_0996_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5704_ (.I(_0996_),
    .Z(_0997_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _5705_ (.A1(_0441_),
    .A2(_0981_),
    .A3(_0982_),
    .ZN(_0998_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_2 _5706_ (.A1(_0997_),
    .A2(_0980_),
    .B1(_0973_),
    .B2(\as2650.r123_2[0][3] ),
    .C(_0998_),
    .ZN(_0999_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5707_ (.I(_0999_),
    .Z(_1000_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5708_ (.A1(\as2650.stack[6][11] ),
    .A2(_0986_),
    .ZN(_1001_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _5709_ (.A1(_0963_),
    .A2(_1000_),
    .B(_1001_),
    .ZN(_0019_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5710_ (.I(\as2650.pc[12] ),
    .Z(_1002_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5711_ (.I(_1002_),
    .Z(_1003_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _5712_ (.A1(_0540_),
    .A2(_4416_),
    .A3(_0982_),
    .ZN(_1004_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_1 _5713_ (.A1(_1003_),
    .A2(_0980_),
    .B1(_0972_),
    .B2(\as2650.r123_2[0][4] ),
    .C(_1004_),
    .ZN(_1005_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5714_ (.I(_1005_),
    .Z(_1006_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5715_ (.A1(\as2650.stack[6][12] ),
    .A2(_0986_),
    .ZN(_1007_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _5716_ (.A1(_0977_),
    .A2(_1006_),
    .B(_1007_),
    .ZN(_0020_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5717_ (.I(\as2650.pc[13] ),
    .Z(_1008_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5718_ (.I(_0971_),
    .Z(_1009_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _5719_ (.A1(_0635_),
    .A2(_4416_),
    .A3(_1009_),
    .ZN(_1010_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_1 _5720_ (.A1(_1008_),
    .A2(_0858_),
    .B1(_0972_),
    .B2(\as2650.r123_2[0][5] ),
    .C(_1010_),
    .ZN(_1011_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5721_ (.I(_1011_),
    .Z(_1012_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5722_ (.A1(\as2650.stack[6][13] ),
    .A2(_0962_),
    .ZN(_1013_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _5723_ (.A1(_0977_),
    .A2(_1012_),
    .B(_1013_),
    .ZN(_0021_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _5724_ (.A1(_0715_),
    .A2(_4416_),
    .A3(_1009_),
    .ZN(_1014_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_1 _5725_ (.A1(\as2650.pc[14] ),
    .A2(_0858_),
    .B1(_0972_),
    .B2(\as2650.r123_2[0][6] ),
    .C(_1014_),
    .ZN(_1015_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5726_ (.I(_1015_),
    .Z(_1016_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5727_ (.A1(\as2650.stack[6][14] ),
    .A2(_0962_),
    .ZN(_1017_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _5728_ (.A1(_0977_),
    .A2(_1016_),
    .B(_1017_),
    .ZN(_0022_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5729_ (.A1(_0866_),
    .A2(_4466_),
    .ZN(_1018_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5730_ (.I(_0959_),
    .Z(_1019_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5731_ (.A1(_1018_),
    .A2(_1019_),
    .ZN(_1020_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5732_ (.I(_1020_),
    .Z(_1021_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5733_ (.I(_1021_),
    .Z(_1022_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5734_ (.I(_1021_),
    .Z(_1023_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5735_ (.A1(\as2650.stack[5][8] ),
    .A2(_1023_),
    .ZN(_1024_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _5736_ (.A1(_0976_),
    .A2(_1022_),
    .B(_1024_),
    .ZN(_0023_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5737_ (.I(_1020_),
    .Z(_1025_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5738_ (.A1(\as2650.stack[5][9] ),
    .A2(_1025_),
    .ZN(_1026_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _5739_ (.A1(_0985_),
    .A2(_1022_),
    .B(_1026_),
    .ZN(_0024_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5740_ (.A1(\as2650.stack[5][10] ),
    .A2(_1025_),
    .ZN(_1027_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _5741_ (.A1(_0993_),
    .A2(_1022_),
    .B(_1027_),
    .ZN(_0025_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5742_ (.A1(\as2650.stack[5][11] ),
    .A2(_1025_),
    .ZN(_1028_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _5743_ (.A1(_1000_),
    .A2(_1022_),
    .B(_1028_),
    .ZN(_0026_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5744_ (.A1(\as2650.stack[5][12] ),
    .A2(_1025_),
    .ZN(_1029_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _5745_ (.A1(_1006_),
    .A2(_1023_),
    .B(_1029_),
    .ZN(_0027_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5746_ (.A1(\as2650.stack[5][13] ),
    .A2(_1021_),
    .ZN(_1030_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _5747_ (.A1(_1012_),
    .A2(_1023_),
    .B(_1030_),
    .ZN(_0028_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5748_ (.A1(\as2650.stack[5][14] ),
    .A2(_1021_),
    .ZN(_1031_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _5749_ (.A1(_1016_),
    .A2(_1023_),
    .B(_1031_),
    .ZN(_0029_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5750_ (.I(\as2650.r123_2[0][0] ),
    .ZN(_1032_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _5751_ (.I(_4150_),
    .Z(_1033_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5752_ (.I(_4200_),
    .Z(_1034_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _5753_ (.A1(_1033_),
    .A2(_1034_),
    .ZN(_1035_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5754_ (.A1(_4248_),
    .A2(_4151_),
    .ZN(_1036_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5755_ (.A1(_4143_),
    .A2(_1036_),
    .ZN(_1037_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5756_ (.A1(_4189_),
    .A2(_1037_),
    .ZN(_1038_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5757_ (.A1(_4407_),
    .A2(_1037_),
    .ZN(_1039_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _5758_ (.A1(_4149_),
    .A2(_4198_),
    .A3(_4151_),
    .ZN(_1040_));
 gf180mcu_fd_sc_mcu7t5v0__or4_1 _5759_ (.A1(_4157_),
    .A2(_4242_),
    .A3(_4245_),
    .A4(_1040_),
    .Z(_1041_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _5760_ (.A1(_4210_),
    .A2(_1040_),
    .ZN(_1042_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5761_ (.A1(_0876_),
    .A2(_0688_),
    .ZN(_1043_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_2 _5762_ (.A1(_4180_),
    .A2(_4249_),
    .A3(_4341_),
    .ZN(_1044_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _5763_ (.A1(_1043_),
    .A2(_1044_),
    .ZN(_1045_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _5764_ (.A1(_4223_),
    .A2(_1045_),
    .ZN(_1046_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _5765_ (.A1(_4150_),
    .A2(_4261_),
    .Z(_1047_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5766_ (.A1(_4195_),
    .A2(_1042_),
    .ZN(_1048_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5767_ (.A1(_1047_),
    .A2(_1048_),
    .ZN(_1049_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _5768_ (.A1(_1042_),
    .A2(_1046_),
    .B(_1049_),
    .ZN(_1050_));
 gf180mcu_fd_sc_mcu7t5v0__and4_1 _5769_ (.A1(_1038_),
    .A2(_1039_),
    .A3(_1041_),
    .A4(_1050_),
    .Z(_1051_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5770_ (.A1(_4137_),
    .A2(_1051_),
    .ZN(_1052_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_2 _5771_ (.A1(_4437_),
    .A2(_1035_),
    .B(_1052_),
    .C(_4438_),
    .ZN(_1053_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5772_ (.I(_1053_),
    .Z(_1054_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5773_ (.I(_1054_),
    .Z(_1055_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5774_ (.I(_1052_),
    .Z(_1056_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5775_ (.I(_1041_),
    .Z(_1057_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5776_ (.I(_1039_),
    .Z(_1058_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5777_ (.I(_1058_),
    .Z(_1059_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5778_ (.I(_1041_),
    .Z(_1060_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5779_ (.I(_1039_),
    .Z(_1061_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5780_ (.I(_1048_),
    .Z(_1062_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5781_ (.I(_1062_),
    .Z(_1063_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5782_ (.I(_4377_),
    .ZN(_1064_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5783_ (.A1(_4220_),
    .A2(_1042_),
    .ZN(_1065_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5784_ (.I(_1065_),
    .Z(_1066_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5785_ (.A1(_4228_),
    .A2(_1042_),
    .ZN(_1067_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5786_ (.I(_1067_),
    .Z(_1068_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5787_ (.I(_1065_),
    .Z(_1069_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5788_ (.A1(_4395_),
    .A2(_1037_),
    .ZN(_1070_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5789_ (.I(_1070_),
    .Z(_1071_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5790_ (.I(_1070_),
    .Z(_1072_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5791_ (.A1(_4398_),
    .A2(_1072_),
    .ZN(_1073_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _5792_ (.A1(_4392_),
    .A2(_1071_),
    .B(_1073_),
    .C(_1067_),
    .ZN(_1074_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _5793_ (.A1(_0301_),
    .A2(_1068_),
    .B(_1069_),
    .C(_1074_),
    .ZN(_1075_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5794_ (.I(_1062_),
    .Z(_1076_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _5795_ (.A1(_1064_),
    .A2(_1066_),
    .B(_1075_),
    .C(_1076_),
    .ZN(_1077_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5796_ (.A1(_4406_),
    .A2(_1063_),
    .B(_1077_),
    .ZN(_1078_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5797_ (.A1(_1061_),
    .A2(_1078_),
    .ZN(_1079_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _5798_ (.A1(_4361_),
    .A2(_1059_),
    .B(_1060_),
    .C(_1079_),
    .ZN(_1080_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5799_ (.A1(_4353_),
    .A2(_1057_),
    .B(_1080_),
    .ZN(_1081_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5800_ (.I(_1047_),
    .Z(_1082_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _5801_ (.I(_1082_),
    .Z(_1083_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _5802_ (.I0(_4344_),
    .I1(_1081_),
    .S(_1083_),
    .Z(_1084_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5803_ (.A1(_4472_),
    .A2(_4484_),
    .ZN(_1085_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5804_ (.I(_4170_),
    .Z(_1086_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5805_ (.A1(_1086_),
    .A2(_0341_),
    .ZN(_1087_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5806_ (.A1(_1087_),
    .A2(_1036_),
    .ZN(_1088_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5807_ (.I(_0294_),
    .Z(_1089_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _5808_ (.A1(_1089_),
    .A2(_0969_),
    .A3(_4492_),
    .ZN(_1090_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _5809_ (.A1(_4295_),
    .A2(_0621_),
    .B1(_1085_),
    .B2(_1088_),
    .C(_1090_),
    .ZN(_1091_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _5810_ (.A1(_1056_),
    .A2(_1084_),
    .B(_1091_),
    .C(_1054_),
    .ZN(_1092_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _5811_ (.A1(_1032_),
    .A2(_1055_),
    .B(_1092_),
    .ZN(_0030_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5812_ (.I(\as2650.r123_2[0][1] ),
    .ZN(_1093_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _5813_ (.A1(_1033_),
    .A2(_4261_),
    .ZN(_1094_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5814_ (.I(_4233_),
    .Z(_1095_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_2 _5815_ (.A1(_1095_),
    .A2(_4268_),
    .A3(_1040_),
    .ZN(_1096_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5816_ (.I(_1096_),
    .Z(_1097_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5817_ (.A1(_4513_),
    .A2(_1097_),
    .ZN(_1098_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5818_ (.I(_1076_),
    .Z(_1099_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5819_ (.I(_4334_),
    .Z(_1100_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5820_ (.I(_1069_),
    .Z(_1101_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5821_ (.I(_1067_),
    .Z(_1102_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5822_ (.I(_1102_),
    .Z(_1103_));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _5823_ (.I(_4529_),
    .ZN(_1104_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5824_ (.I(_1072_),
    .Z(_1105_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _5825_ (.A1(_0301_),
    .A2(_4534_),
    .Z(_1106_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5826_ (.A1(_1106_),
    .A2(_1071_),
    .ZN(_1107_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _5827_ (.A1(_1104_),
    .A2(_1105_),
    .B(_1107_),
    .C(_1068_),
    .ZN(_1108_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _5828_ (.A1(_0400_),
    .A2(_1103_),
    .B(_1066_),
    .C(_1108_),
    .ZN(_1109_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5829_ (.I(_1062_),
    .Z(_1110_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _5830_ (.A1(_1100_),
    .A2(_1101_),
    .B(_1109_),
    .C(_1110_),
    .ZN(_1111_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _5831_ (.A1(_4542_),
    .A2(_1099_),
    .B(_1111_),
    .C(_1059_),
    .ZN(_1112_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _5832_ (.A1(_1060_),
    .A2(_1098_),
    .A3(_1112_),
    .ZN(_1113_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5833_ (.A1(_0292_),
    .A2(_1057_),
    .B(_1113_),
    .ZN(_1114_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5834_ (.A1(_0321_),
    .A2(_1094_),
    .ZN(_1115_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _5835_ (.A1(_1094_),
    .A2(_1114_),
    .B(_1115_),
    .ZN(_1116_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5836_ (.I(_1090_),
    .Z(_1117_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _5837_ (.I(_0969_),
    .Z(_1118_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _5838_ (.A1(_1089_),
    .A2(_1118_),
    .A3(_4444_),
    .ZN(_1119_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5839_ (.A1(_0335_),
    .A2(_1119_),
    .ZN(_1120_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _5840_ (.A1(_0344_),
    .A2(_1117_),
    .A3(_1120_),
    .ZN(_1121_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _5841_ (.A1(_1056_),
    .A2(_1116_),
    .B(_1121_),
    .C(_1054_),
    .ZN(_1122_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _5842_ (.A1(_1093_),
    .A2(_1055_),
    .B(_1122_),
    .ZN(_0031_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5843_ (.I(\as2650.r123_2[0][2] ),
    .ZN(_1123_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5844_ (.I(_1053_),
    .Z(_1124_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _5845_ (.A1(_0436_),
    .A2(_1088_),
    .B(_1090_),
    .C(_0437_),
    .ZN(_1125_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5846_ (.I(_1052_),
    .ZN(_1126_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5847_ (.I(_1065_),
    .Z(_1127_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5848_ (.A1(_0378_),
    .A2(_1071_),
    .ZN(_1128_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _5849_ (.A1(_0376_),
    .A2(_1105_),
    .B(_1128_),
    .C(_1102_),
    .ZN(_1129_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _5850_ (.A1(_0372_),
    .A2(_1103_),
    .B(_1127_),
    .C(_1129_),
    .ZN(_1130_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _5851_ (.A1(_4388_),
    .A2(_1101_),
    .B(_1130_),
    .C(_1110_),
    .ZN(_1131_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _5852_ (.A1(_0360_),
    .A2(_1099_),
    .B(_1131_),
    .C(_1061_),
    .ZN(_1132_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5853_ (.A1(_4552_),
    .A2(_1037_),
    .ZN(_1133_));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _5854_ (.I(_1133_),
    .ZN(_1134_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _5855_ (.A1(_0389_),
    .A2(_1097_),
    .B(_1134_),
    .ZN(_1135_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5856_ (.I(_1041_),
    .Z(_1136_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5857_ (.A1(_0358_),
    .A2(_1136_),
    .ZN(_1137_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _5858_ (.A1(_1132_),
    .A2(_1135_),
    .B(_1137_),
    .C(_1094_),
    .ZN(_1138_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _5859_ (.A1(_0422_),
    .A2(_1094_),
    .B(_1138_),
    .ZN(_1139_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5860_ (.A1(_1126_),
    .A2(_1139_),
    .ZN(_1140_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _5861_ (.A1(_1124_),
    .A2(_1125_),
    .A3(_1140_),
    .ZN(_1141_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _5862_ (.A1(_1123_),
    .A2(_1055_),
    .B(_1141_),
    .ZN(_0032_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5863_ (.I(\as2650.r123_2[0][3] ),
    .ZN(_1142_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5864_ (.A1(_0533_),
    .A2(_1119_),
    .ZN(_1143_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _5865_ (.A1(_0536_),
    .A2(_1117_),
    .A3(_1143_),
    .ZN(_1144_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5866_ (.I(_1082_),
    .Z(_1145_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _5867_ (.A1(_4188_),
    .A2(_1040_),
    .ZN(_1146_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5868_ (.I(_0508_),
    .Z(_1147_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5869_ (.A1(_1147_),
    .A2(_1146_),
    .ZN(_1148_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _5870_ (.A1(_0512_),
    .A2(_1146_),
    .B(_1148_),
    .C(_1102_),
    .ZN(_1149_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _5871_ (.A1(_0566_),
    .A2(_1103_),
    .B(_1127_),
    .C(_1149_),
    .ZN(_1150_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _5872_ (.A1(_4527_),
    .A2(_1101_),
    .B(_1150_),
    .C(_1110_),
    .ZN(_1151_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _5873_ (.A1(_0535_),
    .A2(_1099_),
    .B(_1151_),
    .C(_1061_),
    .ZN(_1152_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _5874_ (.A1(_0491_),
    .A2(_1097_),
    .B(_1134_),
    .ZN(_1153_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _5875_ (.A1(_0485_),
    .A2(_1134_),
    .B1(_1152_),
    .B2(_1153_),
    .ZN(_1154_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _5876_ (.A1(_0446_),
    .A2(_0474_),
    .B(_1082_),
    .ZN(_1155_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _5877_ (.A1(_1145_),
    .A2(_1154_),
    .B(_1155_),
    .ZN(_1156_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5878_ (.A1(_1126_),
    .A2(_1156_),
    .ZN(_1157_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _5879_ (.A1(_1124_),
    .A2(_1144_),
    .A3(_1157_),
    .ZN(_1158_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _5880_ (.A1(_1142_),
    .A2(_1055_),
    .B(_1158_),
    .ZN(_0033_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5881_ (.I(\as2650.r123_2[0][4] ),
    .ZN(_1159_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5882_ (.I(_1054_),
    .Z(_1160_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _5883_ (.A1(_0617_),
    .A2(_0621_),
    .B1(_0632_),
    .B2(_1088_),
    .C(_1090_),
    .ZN(_1161_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5884_ (.A1(_0603_),
    .A2(_1070_),
    .ZN(_1162_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5885_ (.I(_4228_),
    .Z(_1163_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_4 _5886_ (.A1(_1033_),
    .A2(_4420_),
    .A3(_4204_),
    .A4(_4211_),
    .ZN(_1164_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5887_ (.A1(_1163_),
    .A2(_1164_),
    .ZN(_1165_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _5888_ (.A1(_0596_),
    .A2(_1072_),
    .B(_1162_),
    .C(_1165_),
    .ZN(_1166_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _5889_ (.A1(_0592_),
    .A2(_1068_),
    .B(_1069_),
    .C(_1166_),
    .ZN(_1167_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5890_ (.A1(_0371_),
    .A2(_1127_),
    .B(_1167_),
    .ZN(_1168_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5891_ (.A1(_1076_),
    .A2(_1168_),
    .ZN(_1169_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _5892_ (.A1(_0500_),
    .A2(_1063_),
    .B(_1169_),
    .C(_1058_),
    .ZN(_1170_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5893_ (.A1(_0578_),
    .A2(_1096_),
    .ZN(_1171_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _5894_ (.A1(_1136_),
    .A2(_1170_),
    .A3(_1171_),
    .ZN(_1172_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5895_ (.A1(_0614_),
    .A2(_1060_),
    .B(_1172_),
    .ZN(_1173_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _5896_ (.I0(_0570_),
    .I1(_1173_),
    .S(_1145_),
    .Z(_1174_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5897_ (.A1(_1126_),
    .A2(_1174_),
    .ZN(_1175_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _5898_ (.A1(_1124_),
    .A2(_1161_),
    .A3(_1175_),
    .ZN(_1176_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _5899_ (.A1(_1159_),
    .A2(_1160_),
    .B(_1176_),
    .ZN(_0034_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5900_ (.I(\as2650.r123_2[0][5] ),
    .ZN(_1177_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5901_ (.A1(_0709_),
    .A2(_1119_),
    .ZN(_1178_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _5902_ (.A1(_0712_),
    .A2(_1117_),
    .A3(_1178_),
    .ZN(_1179_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5903_ (.I(_0683_),
    .Z(_1180_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5904_ (.A1(_1180_),
    .A2(_1146_),
    .ZN(_1181_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _5905_ (.A1(_0690_),
    .A2(_1146_),
    .B(_1181_),
    .C(_1102_),
    .ZN(_1182_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _5906_ (.A1(_0718_),
    .A2(_1068_),
    .B(_1069_),
    .C(_1182_),
    .ZN(_1183_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _5907_ (.A1(_0505_),
    .A2(_1066_),
    .B(_1183_),
    .C(_1076_),
    .ZN(_1184_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _5908_ (.A1(_0670_),
    .A2(_1063_),
    .B(_1184_),
    .C(_1058_),
    .ZN(_1185_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5909_ (.A1(_0698_),
    .A2(_1096_),
    .ZN(_1186_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _5910_ (.A1(_1136_),
    .A2(_1185_),
    .A3(_1186_),
    .ZN(_1187_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5911_ (.A1(_0668_),
    .A2(_1060_),
    .B(_1187_),
    .ZN(_1188_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _5912_ (.I0(_0662_),
    .I1(_1188_),
    .S(_1082_),
    .Z(_1189_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5913_ (.A1(_1126_),
    .A2(_1189_),
    .ZN(_1190_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _5914_ (.A1(_1124_),
    .A2(_1179_),
    .A3(_1190_),
    .ZN(_1191_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _5915_ (.A1(_1177_),
    .A2(_1160_),
    .B(_1191_),
    .ZN(_0035_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5916_ (.I(\as2650.r123_2[0][6] ),
    .ZN(_1192_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5917_ (.A1(_0763_),
    .A2(_1105_),
    .ZN(_1193_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _5918_ (.A1(_0759_),
    .A2(_1105_),
    .B(_1193_),
    .C(_1165_),
    .ZN(_1194_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _5919_ (.A1(_0753_),
    .A2(_1103_),
    .B(_1066_),
    .C(_1194_),
    .ZN(_1195_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5920_ (.A1(_0639_),
    .A2(_1101_),
    .B(_1195_),
    .ZN(_1196_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5921_ (.A1(_0751_),
    .A2(_1063_),
    .B(_1061_),
    .ZN(_1197_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _5922_ (.A1(_1099_),
    .A2(_1196_),
    .B(_1197_),
    .ZN(_1198_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_2 _5923_ (.A1(_0771_),
    .A2(_1097_),
    .B(_1134_),
    .C(_1198_),
    .ZN(_1199_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5924_ (.A1(_0749_),
    .A2(_1057_),
    .B(_1145_),
    .ZN(_1200_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_2 _5925_ (.A1(_0740_),
    .A2(_1083_),
    .B1(_1199_),
    .B2(_1200_),
    .ZN(_1201_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5926_ (.A1(_0781_),
    .A2(_1119_),
    .ZN(_1202_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _5927_ (.A1(_0783_),
    .A2(_1117_),
    .A3(_1202_),
    .ZN(_1203_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _5928_ (.A1(_1056_),
    .A2(_1201_),
    .B(_1203_),
    .C(_1053_),
    .ZN(_1204_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _5929_ (.A1(_1192_),
    .A2(_1160_),
    .B(_1204_),
    .ZN(_0036_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5930_ (.I(\as2650.r123_2[0][7] ),
    .ZN(_1205_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _5931_ (.A1(_0724_),
    .A2(_0797_),
    .B(_0794_),
    .ZN(_1206_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _5932_ (.A1(_0796_),
    .A2(_0800_),
    .A3(_0798_),
    .ZN(_1207_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5933_ (.A1(_1206_),
    .A2(_1207_),
    .B(_0555_),
    .ZN(_1208_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _5934_ (.A1(_0544_),
    .A2(_0807_),
    .B(_0812_),
    .ZN(_1209_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_2 _5935_ (.A1(_1208_),
    .A2(_1209_),
    .B1(_0815_),
    .B2(_0651_),
    .ZN(_1210_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5936_ (.A1(_0473_),
    .A2(_0819_),
    .ZN(_1211_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_4 _5937_ (.A1(_0473_),
    .A2(_0801_),
    .B1(_1210_),
    .B2(_1211_),
    .ZN(_1212_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5938_ (.A1(_0836_),
    .A2(_1072_),
    .B(_1067_),
    .ZN(_1213_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _5939_ (.A1(_0834_),
    .A2(_1071_),
    .B(_1213_),
    .ZN(_1214_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5940_ (.A1(_0516_),
    .A2(_1164_),
    .ZN(_1215_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5941_ (.A1(_0840_),
    .A2(_1165_),
    .B(_1215_),
    .ZN(_1216_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_1 _5942_ (.A1(_0680_),
    .A2(_1127_),
    .B1(_1214_),
    .B2(_1216_),
    .C(_1062_),
    .ZN(_1217_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5943_ (.A1(_0789_),
    .A2(_1110_),
    .B(_1217_),
    .ZN(_1218_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5944_ (.A1(_1058_),
    .A2(_1218_),
    .ZN(_1219_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _5945_ (.A1(_0830_),
    .A2(_1059_),
    .B(_1136_),
    .C(_1219_),
    .ZN(_1220_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5946_ (.A1(_0828_),
    .A2(_1057_),
    .B(_1220_),
    .ZN(_1221_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5947_ (.A1(_1083_),
    .A2(_1221_),
    .ZN(_1222_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _5948_ (.A1(_1212_),
    .A2(_1083_),
    .B(_1222_),
    .ZN(_1223_));
 gf180mcu_fd_sc_mcu7t5v0__and4_1 _5949_ (.A1(_1089_),
    .A2(_1118_),
    .A3(_4492_),
    .A4(_0792_),
    .Z(_1224_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _5950_ (.A1(_1056_),
    .A2(_1223_),
    .B(_1224_),
    .C(_1053_),
    .ZN(_1225_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _5951_ (.A1(_1205_),
    .A2(_1160_),
    .B(_1225_),
    .ZN(_0037_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5952_ (.I(\as2650.psu[5] ),
    .ZN(_1226_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _5953_ (.A1(_0876_),
    .A2(_4157_),
    .A3(_4278_),
    .ZN(_1227_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5954_ (.I(_1227_),
    .Z(_1228_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5955_ (.I(_1228_),
    .Z(_1229_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _5956_ (.I(_4185_),
    .Z(_1230_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _5957_ (.A1(_4219_),
    .A2(_4227_),
    .ZN(_1231_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5958_ (.A1(_1230_),
    .A2(_1231_),
    .ZN(_1232_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5959_ (.I(_1232_),
    .Z(_1233_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5960_ (.I(_4443_),
    .Z(_1234_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5961_ (.I(_4433_),
    .Z(_1235_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _5962_ (.A1(_4426_),
    .A2(_1235_),
    .A3(_4489_),
    .ZN(_1236_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _5963_ (.I(_0854_),
    .Z(_1237_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5964_ (.I(_4197_),
    .Z(_1238_));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _5965_ (.I(_4136_),
    .ZN(_1239_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5966_ (.A1(_1238_),
    .A2(_1239_),
    .ZN(_1240_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _5967_ (.A1(_0469_),
    .A2(_1240_),
    .A3(_4432_),
    .ZN(_1241_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5968_ (.I(_4427_),
    .Z(_1242_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _5969_ (.A1(_4137_),
    .A2(_1242_),
    .A3(_4425_),
    .ZN(_1243_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _5970_ (.A1(_1237_),
    .A2(_1241_),
    .A3(_1243_),
    .ZN(_1244_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _5971_ (.A1(_1234_),
    .A2(_1236_),
    .A3(_1244_),
    .ZN(_1245_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _5972_ (.A1(_1229_),
    .A2(_1233_),
    .A3(_1245_),
    .ZN(_1246_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5973_ (.A1(_0868_),
    .A2(_4423_),
    .ZN(_1247_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5974_ (.I(_1247_),
    .Z(_1248_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5975_ (.I(_1248_),
    .Z(_1249_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5976_ (.I(_4417_),
    .Z(_1250_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5977_ (.I(_1250_),
    .Z(_1251_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5978_ (.I(_1251_),
    .Z(_1252_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5979_ (.A1(_1238_),
    .A2(_4136_),
    .ZN(_1253_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _5980_ (.A1(\as2650.psl[6] ),
    .A2(_4428_),
    .Z(_1254_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _5981_ (.A1(\as2650.psl[7] ),
    .A2(_1239_),
    .Z(_1255_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _5982_ (.A1(_1254_),
    .A2(_1255_),
    .ZN(_1256_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5983_ (.A1(_1253_),
    .A2(_1256_),
    .ZN(_1257_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _5984_ (.A1(_0814_),
    .A2(_1252_),
    .A3(_1257_),
    .ZN(_1258_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5985_ (.A1(_1249_),
    .A2(_1258_),
    .ZN(_1259_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5986_ (.I(_4393_),
    .Z(_1260_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5987_ (.I(_4369_),
    .Z(_1261_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5988_ (.A1(_4215_),
    .A2(_4223_),
    .ZN(_1262_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _5989_ (.A1(_0874_),
    .A2(_4330_),
    .A3(_1262_),
    .ZN(_1263_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5990_ (.I(_1263_),
    .Z(_1264_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _5991_ (.A1(_1261_),
    .A2(_1264_),
    .B(_1233_),
    .C(_1228_),
    .ZN(_1265_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _5992_ (.A1(_1260_),
    .A2(_1265_),
    .Z(_1266_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _5993_ (.A1(_4174_),
    .A2(_4167_),
    .ZN(_1267_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _5994_ (.I(_1267_),
    .Z(_1268_));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _5995_ (.I(_1236_),
    .ZN(_1269_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_4 _5996_ (.A1(_4201_),
    .A2(_1268_),
    .A3(_1269_),
    .A4(_1237_),
    .ZN(_1270_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _5997_ (.I(_4543_),
    .Z(_1271_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5998_ (.I(_1271_),
    .Z(_1272_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5999_ (.I(_1243_),
    .Z(_1273_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _6000_ (.A1(_1272_),
    .A2(_1273_),
    .ZN(_1274_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _6001_ (.I(_0879_),
    .Z(_1275_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _6002_ (.I(_1275_),
    .Z(_1276_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _6003_ (.I(_1276_),
    .Z(_1277_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6004_ (.I(_0874_),
    .Z(_1278_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6005_ (.I(_1262_),
    .Z(_1279_));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _6006_ (.A1(_1278_),
    .A2(_0418_),
    .A3(_1279_),
    .Z(_1280_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6007_ (.A1(_4430_),
    .A2(_1280_),
    .ZN(_1281_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6008_ (.A1(_4214_),
    .A2(_4250_),
    .ZN(_1282_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _6009_ (.I(_1282_),
    .Z(_1283_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _6010_ (.A1(_1277_),
    .A2(_1281_),
    .B(_1233_),
    .C(_1283_),
    .ZN(_1284_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _6011_ (.A1(_1270_),
    .A2(_1274_),
    .A3(_1284_),
    .ZN(_1285_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_2 _6012_ (.A1(_1246_),
    .A2(_1259_),
    .A3(_1266_),
    .A4(_1285_),
    .ZN(_1286_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6013_ (.I(_1229_),
    .Z(_1287_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6014_ (.I(_1086_),
    .Z(_1288_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6015_ (.I(_1288_),
    .Z(_1289_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6016_ (.A1(_0670_),
    .A2(_1289_),
    .ZN(_1290_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6017_ (.I(_0685_),
    .Z(_1291_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _6018_ (.I(_1291_),
    .Z(_1292_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _6019_ (.I(_4443_),
    .Z(_1293_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _6020_ (.I(_1293_),
    .Z(_1294_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _6021_ (.I(_1294_),
    .Z(_1295_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6022_ (.A1(_4199_),
    .A2(_1264_),
    .ZN(_1296_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6023_ (.A1(_1291_),
    .A2(_1296_),
    .ZN(_1297_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _6024_ (.A1(\as2650.psu[5] ),
    .A2(_1292_),
    .B(_1295_),
    .C(_1297_),
    .ZN(_1298_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6025_ (.A1(_1290_),
    .A2(_1298_),
    .ZN(_1299_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _6026_ (.A1(_1287_),
    .A2(_1299_),
    .B(_1286_),
    .ZN(_1300_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6027_ (.I(_4438_),
    .Z(_1301_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _6028_ (.I(_1301_),
    .Z(_1302_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _6029_ (.A1(_1226_),
    .A2(_1286_),
    .B(_1300_),
    .C(_1302_),
    .ZN(_0038_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _6030_ (.I(\as2650.cycle[7] ),
    .Z(_1303_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _6031_ (.I(_4166_),
    .Z(_1304_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _6032_ (.I(_4252_),
    .Z(_1305_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_2 _6033_ (.A1(_4238_),
    .A2(_0886_),
    .A3(_1304_),
    .A4(_1305_),
    .ZN(_1306_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6034_ (.A1(_1303_),
    .A2(_1306_),
    .ZN(_1307_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6035_ (.A1(_4263_),
    .A2(_1307_),
    .ZN(_1308_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _6036_ (.I(_0888_),
    .Z(_1309_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6037_ (.A1(_4254_),
    .A2(_0878_),
    .ZN(_1310_));
 gf180mcu_fd_sc_mcu7t5v0__and4_1 _6038_ (.A1(_1303_),
    .A2(_0886_),
    .A3(_1304_),
    .A4(_1305_),
    .Z(_1311_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_2 _6039_ (.A1(_1309_),
    .A2(_1310_),
    .A3(_1311_),
    .ZN(_1312_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6040_ (.A1(_1308_),
    .A2(_1312_),
    .ZN(_1313_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _6041_ (.A1(_4235_),
    .A2(_4241_),
    .B(_1313_),
    .ZN(_1314_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _6042_ (.I(_4232_),
    .Z(_1315_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _6043_ (.I(_1315_),
    .Z(_1316_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _6044_ (.A1(_1316_),
    .A2(_1267_),
    .ZN(_1317_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6045_ (.A1(_1314_),
    .A2(_1317_),
    .ZN(_1318_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _6046_ (.I(_1034_),
    .Z(_1319_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _6047_ (.I(_4214_),
    .Z(_1320_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _6048_ (.A1(_1320_),
    .A2(_1228_),
    .ZN(_1321_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6049_ (.I(_1315_),
    .Z(_1322_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6050_ (.I(_1322_),
    .Z(_1323_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _6051_ (.I(_0889_),
    .Z(_1324_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6052_ (.A1(_4174_),
    .A2(_4207_),
    .ZN(_1325_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6053_ (.A1(_0883_),
    .A2(_1325_),
    .ZN(_1326_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _6054_ (.I(_1326_),
    .Z(_1327_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6055_ (.A1(_1316_),
    .A2(_1327_),
    .ZN(_1328_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _6056_ (.I(_4235_),
    .Z(_1329_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6057_ (.A1(_1329_),
    .A2(_1306_),
    .ZN(_1330_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6058_ (.A1(_1328_),
    .A2(_1330_),
    .ZN(_1331_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6059_ (.A1(_1323_),
    .A2(_1324_),
    .B(_1331_),
    .ZN(_1332_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_2 _6060_ (.A1(_1319_),
    .A2(_1321_),
    .A3(_1332_),
    .ZN(_1333_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6061_ (.A1(_1318_),
    .A2(_1333_),
    .ZN(_1334_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6062_ (.I(net3),
    .Z(_1335_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _6063_ (.I(_1335_),
    .Z(_1336_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_4 _6064_ (.A1(_1303_),
    .A2(_0886_),
    .A3(_1304_),
    .A4(_1305_),
    .ZN(_1337_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6065_ (.A1(_4238_),
    .A2(_1337_),
    .ZN(_1338_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6066_ (.A1(_1336_),
    .A2(_1338_),
    .ZN(_1339_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _6067_ (.I(_0881_),
    .Z(_1340_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6068_ (.I(_4263_),
    .Z(_1341_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6069_ (.A1(_1340_),
    .A2(_1341_),
    .ZN(_1342_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _6070_ (.A1(_1339_),
    .A2(_1342_),
    .B(_1323_),
    .ZN(_1343_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6071_ (.A1(_1322_),
    .A2(_1086_),
    .ZN(_1344_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6072_ (.A1(_1307_),
    .A2(_1344_),
    .ZN(_1345_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _6073_ (.I(_4167_),
    .Z(_1346_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _6074_ (.A1(_1346_),
    .A2(_4237_),
    .ZN(_1347_));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _6075_ (.I(_4164_),
    .ZN(_1348_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_4 _6076_ (.A1(\as2650.cycle[3] ),
    .A2(_1348_),
    .A3(_4174_),
    .A4(_4172_),
    .ZN(_1349_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_2 _6077_ (.A1(_0883_),
    .A2(_1315_),
    .A3(_1349_),
    .ZN(_1350_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6078_ (.A1(_1347_),
    .A2(_1350_),
    .ZN(_1351_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6079_ (.A1(_1345_),
    .A2(_1351_),
    .ZN(_1352_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _6080_ (.A1(_1343_),
    .A2(_1352_),
    .Z(_1353_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _6081_ (.I(_4168_),
    .Z(_1354_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _6082_ (.I(_4207_),
    .Z(_1355_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _6083_ (.I(_1355_),
    .Z(_1356_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _6084_ (.A1(_1355_),
    .A2(_1305_),
    .ZN(_1357_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6085_ (.A1(_4551_),
    .A2(_1357_),
    .ZN(_1358_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _6086_ (.A1(_1354_),
    .A2(_1356_),
    .A3(_1358_),
    .ZN(_1359_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6087_ (.A1(_4215_),
    .A2(_0874_),
    .ZN(_1360_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6088_ (.A1(_1360_),
    .A2(_1227_),
    .ZN(_1361_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6089_ (.A1(_4394_),
    .A2(_1361_),
    .ZN(_1362_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6090_ (.A1(_4550_),
    .A2(_0879_),
    .ZN(_1363_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _6091_ (.A1(_1315_),
    .A2(_0882_),
    .ZN(_1364_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _6092_ (.A1(_1282_),
    .A2(_1362_),
    .B(_1363_),
    .C(_1364_),
    .ZN(_1365_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6093_ (.A1(_1359_),
    .A2(_1365_),
    .ZN(_1366_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _6094_ (.I(_4194_),
    .Z(_1367_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _6095_ (.A1(_4442_),
    .A2(_1228_),
    .ZN(_1368_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6096_ (.A1(_4328_),
    .A2(_1230_),
    .ZN(_1369_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _6097_ (.I(_1369_),
    .Z(_1370_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_2 _6098_ (.A1(_1367_),
    .A2(_1283_),
    .B1(_1368_),
    .B2(_1370_),
    .ZN(_1371_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_4 _6099_ (.A1(_1334_),
    .A2(_1353_),
    .A3(_1366_),
    .A4(_1371_),
    .ZN(_1372_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6100_ (.I(_1372_),
    .Z(_1373_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6101_ (.I(_1323_),
    .Z(_1374_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _6102_ (.A1(_1374_),
    .A2(_4266_),
    .Z(_1375_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6103_ (.I(_1375_),
    .Z(_1376_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6104_ (.I(_1375_),
    .Z(_1377_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6105_ (.A1(_1377_),
    .A2(_1100_),
    .ZN(_1378_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6106_ (.A1(_4441_),
    .A2(_1376_),
    .B(_1378_),
    .ZN(_1379_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6107_ (.I(_1372_),
    .Z(_1380_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6108_ (.A1(net41),
    .A2(_1380_),
    .ZN(_1381_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _6109_ (.A1(_1373_),
    .A2(_1379_),
    .B(_1381_),
    .C(_1302_),
    .ZN(_0039_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _6110_ (.I(_0337_),
    .Z(_1382_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6111_ (.I(_4387_),
    .Z(_1383_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6112_ (.A1(_1377_),
    .A2(_1383_),
    .ZN(_1384_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6113_ (.A1(_1382_),
    .A2(_1376_),
    .B(_1384_),
    .ZN(_1385_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6114_ (.A1(net42),
    .A2(_1380_),
    .ZN(_1386_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _6115_ (.A1(_1373_),
    .A2(_1385_),
    .B(_1386_),
    .C(_1302_),
    .ZN(_0040_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6116_ (.A1(_1377_),
    .A2(_4527_),
    .ZN(_1387_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6117_ (.A1(_0917_),
    .A2(_1376_),
    .B(_1387_),
    .ZN(_1388_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6118_ (.A1(net43),
    .A2(_1380_),
    .ZN(_1389_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6119_ (.I(_4202_),
    .Z(_1390_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6120_ (.I(_1390_),
    .Z(_1391_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6121_ (.I(_1391_),
    .Z(_1392_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _6122_ (.A1(_1373_),
    .A2(_1388_),
    .B(_1389_),
    .C(_1392_),
    .ZN(_0041_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _6123_ (.I(_0464_),
    .Z(_1393_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6124_ (.A1(_1377_),
    .A2(_1393_),
    .ZN(_1394_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6125_ (.A1(_0924_),
    .A2(_1376_),
    .B(_1394_),
    .ZN(_1395_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6126_ (.A1(net44),
    .A2(_1380_),
    .ZN(_1396_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _6127_ (.A1(_1373_),
    .A2(_1395_),
    .B(_1396_),
    .C(_1392_),
    .ZN(_0042_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6128_ (.I(_1372_),
    .Z(_1397_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6129_ (.I(_1375_),
    .Z(_1398_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6130_ (.I(_1375_),
    .Z(_1399_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6131_ (.A1(_1399_),
    .A2(_0694_),
    .ZN(_1400_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6132_ (.A1(_0579_),
    .A2(_1398_),
    .B(_1400_),
    .ZN(_1401_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6133_ (.I(_1372_),
    .Z(_1402_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6134_ (.A1(net45),
    .A2(_1402_),
    .ZN(_1403_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _6135_ (.A1(_1397_),
    .A2(_1401_),
    .B(_1403_),
    .C(_1392_),
    .ZN(_0043_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6136_ (.A1(_1399_),
    .A2(_0593_),
    .ZN(_1404_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6137_ (.A1(_0711_),
    .A2(_1398_),
    .B(_1404_),
    .ZN(_1405_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6138_ (.A1(net19),
    .A2(_1402_),
    .ZN(_1406_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _6139_ (.A1(_1397_),
    .A2(_1405_),
    .B(_1406_),
    .C(_1392_),
    .ZN(_0044_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6140_ (.A1(_1399_),
    .A2(_0681_),
    .ZN(_1407_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6141_ (.A1(_0944_),
    .A2(_1398_),
    .B(_1407_),
    .ZN(_1408_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6142_ (.A1(net20),
    .A2(_1402_),
    .ZN(_1409_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6143_ (.I(_1391_),
    .Z(_1410_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _6144_ (.A1(_1397_),
    .A2(_1408_),
    .B(_1409_),
    .C(_1410_),
    .ZN(_0045_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _6145_ (.I(_0790_),
    .Z(_1411_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6146_ (.A1(_1399_),
    .A2(_0754_),
    .ZN(_1412_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6147_ (.A1(_1411_),
    .A2(_1398_),
    .B(_1412_),
    .ZN(_1413_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6148_ (.A1(net21),
    .A2(_1402_),
    .ZN(_1414_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _6149_ (.A1(_1397_),
    .A2(_1413_),
    .B(_1414_),
    .C(_1410_),
    .ZN(_0046_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6150_ (.A1(_0622_),
    .A2(_1019_),
    .ZN(_1415_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6151_ (.I(_1415_),
    .Z(_1416_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6152_ (.I(_1416_),
    .Z(_1417_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6153_ (.I(_1416_),
    .Z(_1418_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6154_ (.A1(\as2650.stack[4][8] ),
    .A2(_1418_),
    .ZN(_1419_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _6155_ (.A1(_0976_),
    .A2(_1417_),
    .B(_1419_),
    .ZN(_0047_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6156_ (.I(_1415_),
    .Z(_1420_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6157_ (.A1(\as2650.stack[4][9] ),
    .A2(_1420_),
    .ZN(_1421_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _6158_ (.A1(_0985_),
    .A2(_1417_),
    .B(_1421_),
    .ZN(_0048_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6159_ (.A1(\as2650.stack[4][10] ),
    .A2(_1420_),
    .ZN(_1422_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _6160_ (.A1(_0993_),
    .A2(_1417_),
    .B(_1422_),
    .ZN(_0049_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6161_ (.A1(\as2650.stack[4][11] ),
    .A2(_1420_),
    .ZN(_1423_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _6162_ (.A1(_1000_),
    .A2(_1417_),
    .B(_1423_),
    .ZN(_0050_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6163_ (.A1(\as2650.stack[4][12] ),
    .A2(_1420_),
    .ZN(_1424_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _6164_ (.A1(_1006_),
    .A2(_1418_),
    .B(_1424_),
    .ZN(_0051_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6165_ (.A1(\as2650.stack[4][13] ),
    .A2(_1416_),
    .ZN(_1425_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _6166_ (.A1(_1012_),
    .A2(_1418_),
    .B(_1425_),
    .ZN(_0052_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6167_ (.A1(\as2650.stack[4][14] ),
    .A2(_1416_),
    .ZN(_1426_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _6168_ (.A1(_1016_),
    .A2(_1418_),
    .B(_1426_),
    .ZN(_0053_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_1 _6169_ (.A1(_4344_),
    .A2(_0321_),
    .A3(_0422_),
    .A4(_0476_),
    .ZN(_1427_));
 gf180mcu_fd_sc_mcu7t5v0__and4_1 _6170_ (.A1(_0569_),
    .A2(_0662_),
    .A3(_0740_),
    .A4(_1427_),
    .Z(_1428_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _6171_ (.I(_0548_),
    .Z(_1429_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6172_ (.A1(_1429_),
    .A2(_0753_),
    .ZN(_1430_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _6173_ (.A1(_0813_),
    .A2(_1429_),
    .B(_1430_),
    .ZN(_1431_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6174_ (.A1(_4303_),
    .A2(_0403_),
    .B(_0404_),
    .ZN(_1432_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _6175_ (.A1(_0449_),
    .A2(_1432_),
    .B(_0452_),
    .ZN(_1433_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _6176_ (.A1(_0442_),
    .A2(_0467_),
    .B1(_1433_),
    .B2(_0445_),
    .ZN(_1434_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _6177_ (.A1(_0567_),
    .A2(_0561_),
    .B1(_1434_),
    .B2(_0556_),
    .ZN(_1435_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6178_ (.A1(_0641_),
    .A2(_1435_),
    .B(_0722_),
    .ZN(_1436_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _6179_ (.A1(_0721_),
    .A2(_0795_),
    .A3(_1436_),
    .ZN(_1437_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6180_ (.A1(_0810_),
    .A2(_1431_),
    .B(_1437_),
    .ZN(_1438_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6181_ (.A1(\as2650.psl[1] ),
    .A2(_0795_),
    .ZN(_1439_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _6182_ (.A1(_0795_),
    .A2(_0798_),
    .B(_1438_),
    .C(_1439_),
    .ZN(_1440_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _6183_ (.A1(_1438_),
    .A2(_1439_),
    .Z(_1441_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6184_ (.I(_1234_),
    .Z(_1442_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _6185_ (.I(_1442_),
    .Z(_1443_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_1 _6186_ (.A1(_4258_),
    .A2(_1440_),
    .A3(_1441_),
    .B(_1443_),
    .ZN(_1444_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_1 _6187_ (.A1(_0408_),
    .A2(_0445_),
    .A3(_0543_),
    .A4(_0641_),
    .ZN(_1445_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_1 _6188_ (.A1(_1252_),
    .A2(_0403_),
    .A3(_0720_),
    .A4(_0801_),
    .ZN(_1446_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _6189_ (.A1(_4311_),
    .A2(_1445_),
    .A3(_1446_),
    .ZN(_1447_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6190_ (.A1(_1444_),
    .A2(_1447_),
    .ZN(_1448_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_1 _6191_ (.A1(_0600_),
    .A2(_0821_),
    .A3(_1428_),
    .B(_1448_),
    .ZN(_1449_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _6192_ (.I(_1374_),
    .Z(_1450_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _6193_ (.I(_1450_),
    .Z(_1451_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6194_ (.A1(_1322_),
    .A2(_0447_),
    .ZN(_1452_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6195_ (.A1(_0394_),
    .A2(_1452_),
    .ZN(_1453_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _6196_ (.A1(_0360_),
    .A2(_4541_),
    .A3(_4405_),
    .ZN(_1454_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_1 _6197_ (.A1(_0751_),
    .A2(_0669_),
    .A3(_0500_),
    .A4(_0492_),
    .ZN(_1455_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _6198_ (.A1(_1454_),
    .A2(_1455_),
    .B(_0789_),
    .ZN(_1456_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _6199_ (.A1(_0394_),
    .A2(_1452_),
    .Z(_1457_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6200_ (.A1(_0754_),
    .A2(_1457_),
    .ZN(_1458_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6201_ (.A1(_0824_),
    .A2(_1458_),
    .ZN(_1459_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _6202_ (.A1(_1453_),
    .A2(_1456_),
    .B(_1459_),
    .C(_1295_),
    .ZN(_1460_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6203_ (.A1(_1451_),
    .A2(_1460_),
    .ZN(_1461_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _6204_ (.I(_4250_),
    .Z(_1462_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _6205_ (.I(_1462_),
    .Z(_1463_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _6206_ (.I(_0884_),
    .Z(_1464_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6207_ (.A1(_1464_),
    .A2(_1355_),
    .ZN(_1465_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6208_ (.A1(_1320_),
    .A2(_1247_),
    .ZN(_1466_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _6209_ (.A1(_1465_),
    .A2(_1232_),
    .A3(_1466_),
    .ZN(_1467_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _6210_ (.A1(_0393_),
    .A2(_4431_),
    .Z(_1468_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _6211_ (.A1(_0340_),
    .A2(_1468_),
    .B(_1429_),
    .ZN(_1469_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _6212_ (.A1(_4543_),
    .A2(_1361_),
    .ZN(_1470_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _6213_ (.A1(_4255_),
    .A2(_4232_),
    .ZN(_1471_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6214_ (.A1(_4433_),
    .A2(_4489_),
    .ZN(_1472_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _6215_ (.A1(_1471_),
    .A2(_0394_),
    .A3(_1472_),
    .ZN(_1473_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _6216_ (.A1(_1045_),
    .A2(_1470_),
    .A3(_1473_),
    .ZN(_1474_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_2 _6217_ (.A1(_1463_),
    .A2(_1467_),
    .B1(_1469_),
    .B2(_1474_),
    .ZN(_1475_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _6218_ (.A1(_1293_),
    .A2(_0516_),
    .A3(_1229_),
    .ZN(_1476_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_2 _6219_ (.A1(_1095_),
    .A2(_1242_),
    .B1(_4544_),
    .B2(_4199_),
    .ZN(_1477_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6220_ (.A1(_4187_),
    .A2(_1477_),
    .B(_4419_),
    .ZN(_1478_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _6221_ (.I(_1465_),
    .Z(_1479_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _6222_ (.I(_1044_),
    .Z(_1480_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _6223_ (.A1(_1320_),
    .A2(_1250_),
    .ZN(_1481_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _6224_ (.I(_0867_),
    .Z(_1482_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _6225_ (.A1(_1482_),
    .A2(_1369_),
    .ZN(_1483_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_4 _6226_ (.A1(_1479_),
    .A2(_4187_),
    .B1(_1480_),
    .B2(_1481_),
    .C(_1483_),
    .ZN(_1484_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _6227_ (.A1(_1476_),
    .A2(_1478_),
    .A3(_1484_),
    .ZN(_1485_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _6228_ (.I(_1034_),
    .Z(_1486_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_4 _6229_ (.A1(_4551_),
    .A2(_1271_),
    .A3(_0397_),
    .A4(_0339_),
    .ZN(_1487_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6230_ (.A1(_1486_),
    .A2(_1487_),
    .ZN(_1488_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6231_ (.I(_0882_),
    .Z(_1489_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6232_ (.I(_1489_),
    .Z(_1490_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6233_ (.A1(_1490_),
    .A2(_1317_),
    .ZN(_1491_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6234_ (.A1(_1269_),
    .A2(_1237_),
    .ZN(_1492_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_2 _6235_ (.A1(_4550_),
    .A2(_4341_),
    .A3(_0338_),
    .B(_4417_),
    .ZN(_1493_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6236_ (.A1(_4544_),
    .A2(_1453_),
    .ZN(_1494_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _6237_ (.A1(_1323_),
    .A2(_1493_),
    .A3(_1494_),
    .ZN(_1495_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _6238_ (.A1(_1316_),
    .A2(_1275_),
    .B(_1357_),
    .ZN(_1496_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6239_ (.I(_4255_),
    .Z(_1497_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6240_ (.I(_1497_),
    .Z(_1498_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6241_ (.A1(_1498_),
    .A2(_1248_),
    .ZN(_1499_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _6242_ (.I(_4208_),
    .Z(_1500_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _6243_ (.A1(_0884_),
    .A2(_4167_),
    .ZN(_1501_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6244_ (.A1(_1500_),
    .A2(_1501_),
    .ZN(_1502_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _6245_ (.A1(_4442_),
    .A2(_1241_),
    .Z(_1503_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6246_ (.A1(_0867_),
    .A2(_4550_),
    .ZN(_1504_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _6247_ (.A1(_1499_),
    .A2(_1502_),
    .A3(_1503_),
    .A4(_1504_),
    .ZN(_1505_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_2 _6248_ (.A1(_1492_),
    .A2(_1495_),
    .A3(_1496_),
    .A4(_1505_),
    .ZN(_1506_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _6249_ (.A1(_1464_),
    .A2(_0883_),
    .ZN(_1507_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _6250_ (.A1(_1346_),
    .A2(_1507_),
    .ZN(_1508_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _6251_ (.I(_1508_),
    .Z(_1509_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6252_ (.A1(_1238_),
    .A2(_1263_),
    .ZN(_1510_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6253_ (.A1(_1509_),
    .A2(_1510_),
    .ZN(_1511_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_2 _6254_ (.A1(_1488_),
    .A2(_1491_),
    .A3(_1506_),
    .A4(_1511_),
    .ZN(_1512_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _6255_ (.I(_1471_),
    .Z(_1513_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_2 _6256_ (.A1(_0814_),
    .A2(_1513_),
    .A3(_1266_),
    .ZN(_1514_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_4 _6257_ (.A1(_1475_),
    .A2(_1485_),
    .A3(_1512_),
    .A4(_1514_),
    .ZN(_1515_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _6258_ (.I(_1095_),
    .Z(_1516_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _6259_ (.I(_1516_),
    .Z(_1517_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6260_ (.I(_1517_),
    .Z(_1518_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6261_ (.I(_1043_),
    .Z(_1519_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6262_ (.I(_1519_),
    .Z(_1520_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6263_ (.A1(_1064_),
    .A2(_0745_),
    .ZN(_1521_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _6264_ (.A1(_1520_),
    .A2(_0681_),
    .A3(_1521_),
    .ZN(_1522_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6265_ (.I(_4428_),
    .Z(_1523_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _6266_ (.I(_1288_),
    .Z(_1524_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6267_ (.I(\as2650.psl[6] ),
    .Z(_1525_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _6268_ (.I(_0758_),
    .Z(_1526_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6269_ (.I(_1280_),
    .Z(_1527_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6270_ (.A1(_1239_),
    .A2(_0759_),
    .ZN(_1528_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _6271_ (.A1(_1525_),
    .A2(_1526_),
    .B(_1527_),
    .C(_1528_),
    .ZN(_1529_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _6272_ (.I(_0751_),
    .ZN(_1530_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6273_ (.A1(_1530_),
    .A2(_1273_),
    .ZN(_1531_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _6274_ (.I(_4418_),
    .Z(_1532_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _6275_ (.A1(_1273_),
    .A2(_1456_),
    .B(_1531_),
    .C(_1532_),
    .ZN(_1533_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_1 _6276_ (.A1(_1523_),
    .A2(_1524_),
    .A3(_1529_),
    .B(_1533_),
    .ZN(_1534_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6277_ (.I(_4227_),
    .Z(_1535_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6278_ (.A1(_1535_),
    .A2(_0840_),
    .ZN(_1536_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6279_ (.I(_0718_),
    .Z(_1537_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6280_ (.A1(_0744_),
    .A2(_1537_),
    .ZN(_1538_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _6281_ (.A1(_1383_),
    .A2(_0754_),
    .A3(_0481_),
    .A4(_1538_),
    .ZN(_1539_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6282_ (.A1(_4328_),
    .A2(_1360_),
    .ZN(_1540_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6283_ (.I(_1540_),
    .Z(_1541_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _6284_ (.A1(_1045_),
    .A2(_1534_),
    .B1(_1536_),
    .B2(_1539_),
    .C(_1541_),
    .ZN(_1542_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6285_ (.A1(_1522_),
    .A2(_1542_),
    .ZN(_1543_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6286_ (.I(_1335_),
    .Z(_1544_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6287_ (.I(_1544_),
    .Z(_1545_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _6288_ (.I(_1545_),
    .Z(_1546_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _6289_ (.I(_1540_),
    .Z(_1547_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6290_ (.A1(_1546_),
    .A2(_1547_),
    .ZN(_1548_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _6291_ (.I(_4391_),
    .Z(_1549_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _6292_ (.I(_1549_),
    .Z(_1550_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _6293_ (.I(_1550_),
    .Z(_1551_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _6294_ (.I(_4531_),
    .Z(_1552_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6295_ (.I(_0373_),
    .Z(_1553_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6296_ (.I(_1553_),
    .Z(_1554_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _6297_ (.I(_1554_),
    .Z(_1555_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _6298_ (.I(_1147_),
    .Z(_1556_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_1 _6299_ (.A1(_1551_),
    .A2(_1552_),
    .A3(_1555_),
    .A4(_1556_),
    .ZN(_1557_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6300_ (.I(_0597_),
    .Z(_1558_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6301_ (.I(_1526_),
    .Z(_1559_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _6302_ (.A1(_1558_),
    .A2(_1291_),
    .A3(_1559_),
    .ZN(_1560_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _6303_ (.A1(_1547_),
    .A2(_1557_),
    .A3(_1560_),
    .ZN(_1561_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _6304_ (.A1(_1518_),
    .A2(_1543_),
    .A3(_1548_),
    .A4(_1561_),
    .ZN(_1562_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6305_ (.A1(_1515_),
    .A2(_1562_),
    .ZN(_1563_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _6306_ (.A1(_1449_),
    .A2(_1461_),
    .B(_1563_),
    .ZN(_1564_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6307_ (.I(_4203_),
    .Z(_1565_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _6308_ (.I(_1565_),
    .Z(_1566_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6309_ (.A1(_1525_),
    .A2(_1515_),
    .B(_1566_),
    .ZN(_1567_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6310_ (.A1(_1564_),
    .A2(_1567_),
    .ZN(_0054_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _6311_ (.A1(_4258_),
    .A2(_1212_),
    .B(_1444_),
    .ZN(_1568_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _6312_ (.I(_1462_),
    .Z(_1569_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _6313_ (.I(_1569_),
    .Z(_1570_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6314_ (.I(_1532_),
    .Z(_1571_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6315_ (.I(_1571_),
    .Z(_1572_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _6316_ (.A1(_1411_),
    .A2(_1457_),
    .B(_1458_),
    .C(_1572_),
    .ZN(_1573_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6317_ (.A1(_1570_),
    .A2(_1573_),
    .ZN(_1574_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _6318_ (.I(_1374_),
    .Z(_1575_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6319_ (.I(_1575_),
    .Z(_1576_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6320_ (.A1(_1541_),
    .A2(_1536_),
    .ZN(_1577_));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _6321_ (.A1(_1278_),
    .A2(_4314_),
    .A3(_1279_),
    .Z(_1578_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6322_ (.I(_0837_),
    .Z(_1579_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _6323_ (.I(_0595_),
    .ZN(_1580_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _6324_ (.I(_1580_),
    .Z(_1581_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _6325_ (.I(_1581_),
    .Z(_1582_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _6326_ (.A1(_4463_),
    .A2(_1104_),
    .B1(_0375_),
    .B2(_0849_),
    .ZN(_1583_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _6327_ (.I(net9),
    .ZN(_1584_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6328_ (.I(_1584_),
    .Z(_1585_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _6329_ (.I(_0755_),
    .Z(_1586_));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _6330_ (.I(_1586_),
    .ZN(_1587_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _6331_ (.I(_1587_),
    .Z(_1588_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _6332_ (.I(_4467_),
    .Z(_1589_));
 gf180mcu_fd_sc_mcu7t5v0__oai222_1 _6333_ (.A1(\as2650.psu[3] ),
    .A2(_1585_),
    .B1(_1588_),
    .B2(net27),
    .C1(_1589_),
    .C2(_4392_),
    .ZN(_1590_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _6334_ (.A1(_1226_),
    .A2(_0684_),
    .B(_1583_),
    .C(_1590_),
    .ZN(_1591_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_1 _6335_ (.A1(\as2650.psu[7] ),
    .A2(_1579_),
    .B1(_1582_),
    .B2(\as2650.psu[4] ),
    .C(_1591_),
    .ZN(_1592_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _6336_ (.A1(_1523_),
    .A2(_1578_),
    .A3(_1592_),
    .ZN(_1593_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _6337_ (.I(_1585_),
    .Z(_1594_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _6338_ (.I(\as2650.psl[5] ),
    .ZN(_1595_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _6339_ (.A1(_4316_),
    .A2(_4391_),
    .B1(_0683_),
    .B2(_1595_),
    .ZN(_1596_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_2 _6340_ (.A1(\as2650.overflow ),
    .A2(_0375_),
    .B1(_1594_),
    .B2(_4320_),
    .C(_1596_),
    .ZN(_1597_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _6341_ (.A1(\as2650.psl[1] ),
    .A2(_1104_),
    .B1(_1588_),
    .B2(_1525_),
    .ZN(_1598_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _6342_ (.I(_0835_),
    .Z(_1599_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _6343_ (.A1(\as2650.psl[7] ),
    .A2(_1599_),
    .B1(_1581_),
    .B2(_4248_),
    .ZN(_1600_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _6344_ (.I(_1238_),
    .Z(_1601_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_1 _6345_ (.A1(_1597_),
    .A2(_1598_),
    .A3(_1600_),
    .B(_1601_),
    .ZN(_1602_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6346_ (.A1(_1578_),
    .A2(_1602_),
    .ZN(_1603_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6347_ (.I(net3),
    .Z(_1604_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _6348_ (.I(_1604_),
    .Z(_1605_));
 gf180mcu_fd_sc_mcu7t5v0__aoi222_1 _6349_ (.A1(_1549_),
    .A2(_4334_),
    .B1(_0592_),
    .B2(_0684_),
    .C1(_0753_),
    .C2(_1605_),
    .ZN(_1606_));
 gf180mcu_fd_sc_mcu7t5v0__aoi222_1 _6350_ (.A1(_4530_),
    .A2(_4387_),
    .B1(_4526_),
    .B2(_1554_),
    .C1(_0680_),
    .C2(_0758_),
    .ZN(_1607_));
 gf180mcu_fd_sc_mcu7t5v0__aoi222_1 _6351_ (.A1(_1147_),
    .A2(_1393_),
    .B1(_0505_),
    .B2(_0597_),
    .C1(_1578_),
    .C2(_1601_),
    .ZN(_1608_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _6352_ (.A1(_1606_),
    .A2(_1607_),
    .A3(_1608_),
    .ZN(_1609_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _6353_ (.A1(_1261_),
    .A2(_1527_),
    .B1(_1603_),
    .B2(_1609_),
    .ZN(_1610_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6354_ (.I(\as2650.psl[7] ),
    .Z(_1611_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _6355_ (.I(_1253_),
    .Z(_1612_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _6356_ (.A1(_1611_),
    .A2(_1612_),
    .A3(_1264_),
    .ZN(_1613_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6357_ (.I(_0837_),
    .Z(_1614_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _6358_ (.A1(_1593_),
    .A2(_1610_),
    .B1(_1613_),
    .B2(_1614_),
    .ZN(_1615_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6359_ (.I(net3),
    .Z(_1616_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _6360_ (.I(_1616_),
    .Z(_1617_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6361_ (.I(_1617_),
    .Z(_1618_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _6362_ (.I(_1618_),
    .Z(_1619_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6363_ (.A1(_1619_),
    .A2(_1281_),
    .ZN(_1620_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _6364_ (.A1(_1281_),
    .A2(_1615_),
    .B1(_1620_),
    .B2(_1611_),
    .ZN(_1621_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6365_ (.I(_1442_),
    .Z(_1622_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6366_ (.I(_4219_),
    .Z(_1623_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6367_ (.I(_1623_),
    .Z(_1624_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6368_ (.A1(_1622_),
    .A2(_1624_),
    .ZN(_1625_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6369_ (.A1(_0790_),
    .A2(_1571_),
    .ZN(_1626_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _6370_ (.I(_1519_),
    .Z(_1627_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6371_ (.I(_1480_),
    .Z(_1628_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _6372_ (.A1(_1520_),
    .A2(_1537_),
    .B(_1628_),
    .ZN(_1629_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_1 _6373_ (.A1(_1621_),
    .A2(_1625_),
    .B1(_1626_),
    .B2(_1627_),
    .C(_1629_),
    .ZN(_1630_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6374_ (.A1(_1577_),
    .A2(_1630_),
    .ZN(_1631_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _6375_ (.A1(_1576_),
    .A2(_1548_),
    .A3(_1631_),
    .ZN(_1632_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6376_ (.A1(_1568_),
    .A2(_1574_),
    .B(_1632_),
    .ZN(_1633_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _6377_ (.I(_1565_),
    .Z(_1634_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _6378_ (.I(_1634_),
    .Z(_1635_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6379_ (.A1(_1611_),
    .A2(_1515_),
    .B(_1635_),
    .ZN(_1636_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _6380_ (.A1(_1515_),
    .A2(_1633_),
    .B(_1636_),
    .ZN(_0055_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6381_ (.A1(_4467_),
    .A2(_4463_),
    .ZN(_1637_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6382_ (.I(_1637_),
    .Z(_1638_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6383_ (.I(_1638_),
    .Z(_1639_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6384_ (.I(_1639_),
    .Z(_1640_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _6385_ (.A1(_0851_),
    .A2(_1640_),
    .A3(_1019_),
    .ZN(_1641_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6386_ (.I(_1641_),
    .Z(_1642_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6387_ (.I(_1642_),
    .Z(_1643_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6388_ (.I(_1642_),
    .Z(_1644_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6389_ (.A1(\as2650.stack[3][8] ),
    .A2(_1644_),
    .ZN(_1645_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _6390_ (.A1(_0976_),
    .A2(_1643_),
    .B(_1645_),
    .ZN(_0056_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6391_ (.I(_1641_),
    .Z(_1646_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6392_ (.A1(\as2650.stack[3][9] ),
    .A2(_1646_),
    .ZN(_1647_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _6393_ (.A1(_0985_),
    .A2(_1643_),
    .B(_1647_),
    .ZN(_0057_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6394_ (.A1(\as2650.stack[3][10] ),
    .A2(_1646_),
    .ZN(_1648_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _6395_ (.A1(_0993_),
    .A2(_1643_),
    .B(_1648_),
    .ZN(_0058_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6396_ (.A1(\as2650.stack[3][11] ),
    .A2(_1646_),
    .ZN(_1649_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _6397_ (.A1(_1000_),
    .A2(_1643_),
    .B(_1649_),
    .ZN(_0059_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6398_ (.A1(\as2650.stack[3][12] ),
    .A2(_1646_),
    .ZN(_1650_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _6399_ (.A1(_1006_),
    .A2(_1644_),
    .B(_1650_),
    .ZN(_0060_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6400_ (.A1(\as2650.stack[3][13] ),
    .A2(_1642_),
    .ZN(_1651_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _6401_ (.A1(_1012_),
    .A2(_1644_),
    .B(_1651_),
    .ZN(_0061_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6402_ (.A1(\as2650.stack[3][14] ),
    .A2(_1642_),
    .ZN(_1652_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _6403_ (.A1(_1016_),
    .A2(_1644_),
    .B(_1652_),
    .ZN(_0062_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6404_ (.I(_0975_),
    .Z(_1653_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6405_ (.A1(_4456_),
    .A2(\as2650.psu[1] ),
    .ZN(_1654_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6406_ (.I(_1654_),
    .Z(_1655_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6407_ (.I(_1655_),
    .Z(_1656_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6408_ (.I(_1656_),
    .Z(_1657_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _6409_ (.A1(_0851_),
    .A2(_1657_),
    .A3(_0960_),
    .ZN(_1658_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6410_ (.I(_1658_),
    .Z(_1659_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6411_ (.I(_1659_),
    .Z(_1660_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6412_ (.I(_1659_),
    .Z(_1661_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6413_ (.A1(\as2650.stack[2][8] ),
    .A2(_1661_),
    .ZN(_1662_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _6414_ (.A1(_1653_),
    .A2(_1660_),
    .B(_1662_),
    .ZN(_0063_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6415_ (.I(_0984_),
    .Z(_1663_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6416_ (.I(_1658_),
    .Z(_1664_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6417_ (.A1(\as2650.stack[2][9] ),
    .A2(_1664_),
    .ZN(_1665_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _6418_ (.A1(_1663_),
    .A2(_1660_),
    .B(_1665_),
    .ZN(_0064_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6419_ (.I(_0992_),
    .Z(_1666_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6420_ (.A1(\as2650.stack[2][10] ),
    .A2(_1664_),
    .ZN(_1667_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _6421_ (.A1(_1666_),
    .A2(_1660_),
    .B(_1667_),
    .ZN(_0065_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6422_ (.I(_0999_),
    .Z(_1668_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6423_ (.A1(\as2650.stack[2][11] ),
    .A2(_1664_),
    .ZN(_1669_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _6424_ (.A1(_1668_),
    .A2(_1660_),
    .B(_1669_),
    .ZN(_0066_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6425_ (.I(_1005_),
    .Z(_1670_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6426_ (.A1(\as2650.stack[2][12] ),
    .A2(_1664_),
    .ZN(_1671_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _6427_ (.A1(_1670_),
    .A2(_1661_),
    .B(_1671_),
    .ZN(_0067_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6428_ (.I(_1011_),
    .Z(_1672_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6429_ (.A1(\as2650.stack[2][13] ),
    .A2(_1659_),
    .ZN(_1673_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _6430_ (.A1(_1672_),
    .A2(_1661_),
    .B(_1673_),
    .ZN(_0068_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6431_ (.I(_1015_),
    .Z(_1674_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6432_ (.A1(\as2650.stack[2][14] ),
    .A2(_1659_),
    .ZN(_1675_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _6433_ (.A1(_1674_),
    .A2(_1661_),
    .B(_1675_),
    .ZN(_0069_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _6434_ (.I(_1500_),
    .Z(_1676_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _6435_ (.I(_1676_),
    .Z(_1677_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _6436_ (.I(_1464_),
    .Z(_1678_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6437_ (.I(_1335_),
    .Z(_1679_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _6438_ (.I(_1679_),
    .Z(_1680_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _6439_ (.A1(_1253_),
    .A2(_4431_),
    .ZN(_1681_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6440_ (.A1(_4223_),
    .A2(_1681_),
    .ZN(_1682_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6441_ (.A1(_0876_),
    .A2(_1682_),
    .ZN(_1683_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _6442_ (.I(_1683_),
    .Z(_1684_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6443_ (.I(_1684_),
    .Z(_1685_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6444_ (.A1(_1680_),
    .A2(_1685_),
    .ZN(_1686_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6445_ (.A1(_1678_),
    .A2(_1686_),
    .ZN(_1687_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_4 _6446_ (.A1(_1677_),
    .A2(_1118_),
    .A3(_1356_),
    .A4(_1687_),
    .ZN(_1688_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _6447_ (.I(_1688_),
    .ZN(_1689_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6448_ (.I(_1689_),
    .Z(_1690_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _6449_ (.I(_1551_),
    .Z(_1691_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _6450_ (.I(_1502_),
    .Z(_1692_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6451_ (.A1(_1691_),
    .A2(_1692_),
    .B(_1690_),
    .ZN(_1693_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6452_ (.A1(_1523_),
    .A2(_1690_),
    .B(_1693_),
    .ZN(_0070_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6453_ (.A1(_1552_),
    .A2(_1692_),
    .B(_1689_),
    .ZN(_1694_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6454_ (.A1(_1239_),
    .A2(_1690_),
    .B(_1694_),
    .ZN(_0071_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6455_ (.I(_0877_),
    .Z(_1695_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _6456_ (.I(_1695_),
    .Z(_1696_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_2 _6457_ (.A1(_1678_),
    .A2(_1354_),
    .A3(_0852_),
    .A4(_1346_),
    .ZN(_1697_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6458_ (.I(_1697_),
    .Z(_1698_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _6459_ (.I(_1554_),
    .Z(_1699_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _6460_ (.A1(_1696_),
    .A2(_1688_),
    .B1(_1698_),
    .B2(_1699_),
    .ZN(_1700_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _6461_ (.I(_1700_),
    .ZN(_0072_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _6462_ (.I(_1504_),
    .Z(_1701_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6463_ (.A1(_1502_),
    .A2(_1701_),
    .ZN(_1702_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6464_ (.A1(_1292_),
    .A2(_1692_),
    .B(_1702_),
    .ZN(_1703_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6465_ (.I(_1697_),
    .Z(_1704_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6466_ (.A1(_0814_),
    .A2(_1704_),
    .ZN(_1705_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _6467_ (.A1(_1690_),
    .A2(_1703_),
    .B(_1705_),
    .ZN(_0073_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _6468_ (.I(_1559_),
    .Z(_1706_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _6469_ (.A1(_4160_),
    .A2(_1688_),
    .B1(_1698_),
    .B2(_1706_),
    .ZN(_1707_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _6470_ (.I(_1707_),
    .ZN(_0074_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _6471_ (.I(_1604_),
    .Z(_1708_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6472_ (.I(_1708_),
    .Z(_1709_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6473_ (.I(_1709_),
    .Z(_1710_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _6474_ (.I(_1710_),
    .Z(_1711_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _6475_ (.A1(_4328_),
    .A2(_1688_),
    .B1(_1704_),
    .B2(_1711_),
    .ZN(_1712_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _6476_ (.I(_1712_),
    .ZN(_0075_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _6477_ (.I(_1084_),
    .ZN(_1713_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _6478_ (.A1(_1601_),
    .A2(_1051_),
    .Z(_1714_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6479_ (.I(_1714_),
    .Z(_1715_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6480_ (.A1(_0853_),
    .A2(_4489_),
    .ZN(_1716_));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _6481_ (.I(_1714_),
    .ZN(_1717_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_2 _6482_ (.A1(_1716_),
    .A2(_1035_),
    .B(_1717_),
    .C(_4202_),
    .ZN(_1718_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6483_ (.I(_1718_),
    .Z(_1719_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _6484_ (.I0(\as2650.r123[0][0] ),
    .I1(\as2650.r123_2[0][0] ),
    .S(_4146_),
    .Z(_1720_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6485_ (.I(_1720_),
    .Z(_1721_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6486_ (.I(_1721_),
    .Z(_1722_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6487_ (.I(_1722_),
    .Z(_1723_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _6488_ (.A1(_4405_),
    .A2(_1723_),
    .Z(_1724_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _6489_ (.A1(_0294_),
    .A2(_4152_),
    .A3(_4419_),
    .A4(_1236_),
    .ZN(_1725_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6490_ (.A1(_1725_),
    .A2(_1718_),
    .ZN(_1726_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6491_ (.I(_1726_),
    .Z(_1727_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _6492_ (.A1(\as2650.r123_2[1][0] ),
    .A2(_1719_),
    .B1(_1724_),
    .B2(_1727_),
    .ZN(_1728_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6493_ (.A1(_1713_),
    .A2(_1715_),
    .B(_1728_),
    .ZN(_0076_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6494_ (.I(_1718_),
    .Z(_1729_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _6495_ (.I0(\as2650.r123[0][1] ),
    .I1(\as2650.r123_2[0][1] ),
    .S(_4145_),
    .Z(_1730_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6496_ (.I(_1730_),
    .Z(_1731_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6497_ (.I(_1731_),
    .Z(_1732_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6498_ (.I(_1732_),
    .Z(_1733_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _6499_ (.A1(_4541_),
    .A2(_1733_),
    .A3(_1724_),
    .ZN(_1734_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _6500_ (.I(_1734_),
    .ZN(_1735_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6501_ (.I(_1723_),
    .Z(_1736_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _6502_ (.A1(_0337_),
    .A2(_1736_),
    .B1(_1733_),
    .B2(_4441_),
    .ZN(_1737_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6503_ (.A1(_1735_),
    .A2(_1737_),
    .ZN(_1738_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _6504_ (.A1(\as2650.r123_2[1][1] ),
    .A2(_1729_),
    .B1(_1727_),
    .B2(_1738_),
    .ZN(_1739_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6505_ (.A1(_1116_),
    .A2(_1717_),
    .ZN(_1740_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6506_ (.A1(_1739_),
    .A2(_1740_),
    .ZN(_0077_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6507_ (.I(_1726_),
    .Z(_1741_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6508_ (.A1(_0359_),
    .A2(_1722_),
    .ZN(_1742_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6509_ (.A1(_4541_),
    .A2(_1733_),
    .ZN(_1743_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _6510_ (.I0(\as2650.r123[0][2] ),
    .I1(\as2650.r123_2[0][2] ),
    .S(\as2650.psl[4] ),
    .Z(_1744_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6511_ (.I(_1744_),
    .Z(_1745_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6512_ (.I(_1745_),
    .Z(_1746_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6513_ (.A1(_4284_),
    .A2(_1746_),
    .ZN(_1747_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6514_ (.I(_1745_),
    .Z(_1748_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6515_ (.I(_1748_),
    .Z(_1749_));
 gf180mcu_fd_sc_mcu7t5v0__and4_1 _6516_ (.A1(_4383_),
    .A2(_4294_),
    .A3(_1732_),
    .A4(_1749_),
    .Z(_1750_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _6517_ (.A1(_1743_),
    .A2(_1747_),
    .B(_1750_),
    .ZN(_1751_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _6518_ (.A1(_1742_),
    .A2(_1751_),
    .Z(_1752_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _6519_ (.A1(_1734_),
    .A2(_1752_),
    .Z(_1753_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _6520_ (.A1(\as2650.r123_2[1][2] ),
    .A2(_1719_),
    .B1(_1741_),
    .B2(_1753_),
    .ZN(_1754_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6521_ (.A1(_1139_),
    .A2(_1715_),
    .B(_1754_),
    .ZN(_0078_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6522_ (.A1(_0364_),
    .A2(_1722_),
    .ZN(_1755_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _6523_ (.A1(_1750_),
    .A2(_1755_),
    .Z(_1756_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6524_ (.I(\as2650.r0[1] ),
    .Z(_1757_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6525_ (.A1(_1757_),
    .A2(_1746_),
    .ZN(_1758_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6526_ (.I(\as2650.r0[2] ),
    .Z(_1759_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6527_ (.A1(_1759_),
    .A2(_1731_),
    .ZN(_1760_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _6528_ (.I0(\as2650.r123[0][3] ),
    .I1(\as2650.r123_2[0][3] ),
    .S(_4144_),
    .Z(_1761_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6529_ (.I(_1761_),
    .Z(_1762_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6530_ (.I(_1762_),
    .Z(_1763_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6531_ (.I(_1763_),
    .Z(_1764_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6532_ (.A1(_4405_),
    .A2(_1764_),
    .ZN(_1765_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _6533_ (.A1(_1758_),
    .A2(_1760_),
    .A3(_1765_),
    .Z(_1766_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _6534_ (.A1(_1756_),
    .A2(_1766_),
    .ZN(_1767_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _6535_ (.A1(_0359_),
    .A2(_1723_),
    .A3(_1751_),
    .ZN(_1768_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _6536_ (.A1(_1734_),
    .A2(_1752_),
    .Z(_1769_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6537_ (.A1(_1768_),
    .A2(_1769_),
    .ZN(_1770_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _6538_ (.A1(_1767_),
    .A2(_1770_),
    .Z(_1771_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _6539_ (.I(_1771_),
    .ZN(_1772_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _6540_ (.A1(\as2650.r123_2[1][3] ),
    .A2(_1719_),
    .B1(_1741_),
    .B2(_1772_),
    .ZN(_1773_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6541_ (.A1(_1156_),
    .A2(_1715_),
    .B(_1773_),
    .ZN(_0079_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6542_ (.A1(_1769_),
    .A2(_1767_),
    .ZN(_1774_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _6543_ (.A1(_1768_),
    .A2(_1767_),
    .Z(_1775_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6544_ (.A1(_1757_),
    .A2(_1763_),
    .ZN(_1776_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6545_ (.A1(_0363_),
    .A2(_1732_),
    .ZN(_1777_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6546_ (.A1(_1759_),
    .A2(_1749_),
    .ZN(_1778_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _6547_ (.A1(_1776_),
    .A2(_1777_),
    .A3(_1778_),
    .Z(_1779_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6548_ (.A1(_4146_),
    .A2(\as2650.r123_2[0][4] ),
    .ZN(_1780_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6549_ (.A1(_4147_),
    .A2(_0540_),
    .B(_1780_),
    .ZN(_1781_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _6550_ (.A1(_4285_),
    .A2(_1781_),
    .Z(_1782_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6551_ (.I(_1762_),
    .Z(_1783_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _6552_ (.A1(_4382_),
    .A2(_1748_),
    .B1(_1783_),
    .B2(_4284_),
    .ZN(_1784_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_2 _6553_ (.A1(_1747_),
    .A2(_1776_),
    .B1(_1784_),
    .B2(_1760_),
    .ZN(_1785_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _6554_ (.A1(_0499_),
    .A2(_1721_),
    .Z(_1786_));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_1 _6555_ (.A1(_1782_),
    .A2(_1785_),
    .A3(_1786_),
    .ZN(_1787_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _6556_ (.A1(_0492_),
    .A2(_1722_),
    .A3(_1750_),
    .ZN(_1788_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6557_ (.A1(_1756_),
    .A2(_1766_),
    .B(_1788_),
    .ZN(_1789_));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_1 _6558_ (.A1(_1779_),
    .A2(_1787_),
    .A3(_1789_),
    .ZN(_1790_));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_1 _6559_ (.A1(_1774_),
    .A2(_1775_),
    .A3(_1790_),
    .ZN(_1791_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _6560_ (.I(_1791_),
    .ZN(_1792_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _6561_ (.A1(\as2650.r123_2[1][4] ),
    .A2(_1719_),
    .B1(_1741_),
    .B2(_1792_),
    .ZN(_1793_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6562_ (.A1(_1174_),
    .A2(_1715_),
    .B(_1793_),
    .ZN(_0080_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _6563_ (.A1(_1725_),
    .A2(_1718_),
    .Z(_1794_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6564_ (.I(_1794_),
    .Z(_1795_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6565_ (.A1(_1775_),
    .A2(_1790_),
    .ZN(_1796_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6566_ (.A1(_1775_),
    .A2(_1790_),
    .ZN(_1797_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _6567_ (.A1(_1774_),
    .A2(_1796_),
    .B(_1797_),
    .ZN(_1798_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _6568_ (.A1(_1779_),
    .A2(_1787_),
    .Z(_1799_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6569_ (.A1(_1799_),
    .A2(_1789_),
    .ZN(_1800_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6570_ (.A1(_1779_),
    .A2(_1787_),
    .ZN(_1801_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _6571_ (.A1(_1785_),
    .A2(_1786_),
    .Z(_1802_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _6572_ (.A1(_1785_),
    .A2(_1786_),
    .Z(_1803_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _6573_ (.A1(_1782_),
    .A2(_1802_),
    .B(_1803_),
    .ZN(_1804_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6574_ (.A1(_4519_),
    .A2(_1783_),
    .ZN(_1805_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6575_ (.A1(_0498_),
    .A2(_1731_),
    .ZN(_1806_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6576_ (.A1(_0363_),
    .A2(_1748_),
    .ZN(_1807_));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_1 _6577_ (.A1(_1805_),
    .A2(_1806_),
    .A3(_1807_),
    .ZN(_1808_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _6578_ (.I0(\as2650.r123[0][5] ),
    .I1(\as2650.r123_2[0][5] ),
    .S(_4144_),
    .Z(_1809_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6579_ (.I(_1809_),
    .Z(_1810_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6580_ (.I(_1810_),
    .Z(_1811_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6581_ (.I(_1811_),
    .Z(_1812_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6582_ (.A1(_4294_),
    .A2(_1812_),
    .ZN(_1813_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _6583_ (.A1(_1808_),
    .A2(_1813_),
    .Z(_1814_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6584_ (.A1(_4383_),
    .A2(_1781_),
    .ZN(_1815_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _6585_ (.A1(_1759_),
    .A2(_1746_),
    .B1(_1783_),
    .B2(_1757_),
    .ZN(_1816_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_2 _6586_ (.A1(_1758_),
    .A2(_1805_),
    .B1(_1816_),
    .B2(_1777_),
    .ZN(_1817_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6587_ (.A1(_0585_),
    .A2(_1721_),
    .ZN(_1818_));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_1 _6588_ (.A1(_1815_),
    .A2(_1817_),
    .A3(_1818_),
    .ZN(_1819_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _6589_ (.A1(_1814_),
    .A2(_1819_),
    .Z(_1820_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _6590_ (.A1(_1801_),
    .A2(_1804_),
    .A3(_1820_),
    .Z(_1821_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _6591_ (.A1(_1800_),
    .A2(_1821_),
    .ZN(_1822_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _6592_ (.A1(_1798_),
    .A2(_1822_),
    .ZN(_1823_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6593_ (.A1(_1795_),
    .A2(_1823_),
    .ZN(_1824_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _6594_ (.A1(\as2650.r123_2[1][5] ),
    .A2(_1729_),
    .B(_1824_),
    .ZN(_1825_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6595_ (.A1(_1189_),
    .A2(_1714_),
    .B(_1825_),
    .ZN(_0081_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _6596_ (.A1(_1800_),
    .A2(_1821_),
    .Z(_1826_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6597_ (.A1(_1798_),
    .A2(_1822_),
    .B(_1826_),
    .ZN(_1827_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6598_ (.A1(_1785_),
    .A2(_1786_),
    .ZN(_1828_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6599_ (.A1(_1782_),
    .A2(_1802_),
    .ZN(_1829_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6600_ (.A1(_1828_),
    .A2(_1829_),
    .ZN(_1830_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _6601_ (.A1(_1801_),
    .A2(_1820_),
    .Z(_1831_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _6602_ (.A1(_1801_),
    .A2(_1820_),
    .Z(_1832_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _6603_ (.A1(_1830_),
    .A2(_1831_),
    .B(_1832_),
    .ZN(_1833_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _6604_ (.A1(_0669_),
    .A2(_1736_),
    .B(_1817_),
    .ZN(_1834_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _6605_ (.A1(_0669_),
    .A2(_1723_),
    .A3(_1817_),
    .ZN(_1835_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6606_ (.A1(_1815_),
    .A2(_1834_),
    .B(_1835_),
    .ZN(_1836_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6607_ (.A1(_1814_),
    .A2(_1819_),
    .ZN(_1837_));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _6608_ (.A1(_4294_),
    .A2(_1812_),
    .A3(_1808_),
    .Z(_1838_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6609_ (.A1(_4382_),
    .A2(_1811_),
    .ZN(_1839_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _6610_ (.I0(\as2650.r123[0][6] ),
    .I1(\as2650.r123_2[0][6] ),
    .S(_4145_),
    .Z(_1840_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6611_ (.I(_1840_),
    .Z(_1841_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6612_ (.A1(\as2650.r0[0] ),
    .A2(_1841_),
    .ZN(_1842_));
 gf180mcu_fd_sc_mcu7t5v0__and4_1 _6613_ (.A1(_4382_),
    .A2(_4284_),
    .A3(_1810_),
    .A4(_1841_),
    .Z(_1843_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _6614_ (.A1(_1839_),
    .A2(_1842_),
    .B(_1843_),
    .ZN(_1844_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6615_ (.A1(\as2650.r0[3] ),
    .A2(_1762_),
    .ZN(_1845_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6616_ (.A1(\as2650.r0[5] ),
    .A2(_1730_),
    .ZN(_1846_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6617_ (.A1(\as2650.r0[4] ),
    .A2(_1745_),
    .ZN(_1847_));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_1 _6618_ (.A1(_1845_),
    .A2(_1846_),
    .A3(_1847_),
    .ZN(_1848_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _6619_ (.A1(_1844_),
    .A2(_1848_),
    .Z(_1849_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6620_ (.A1(_4520_),
    .A2(_1781_),
    .ZN(_1850_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _6621_ (.A1(_0363_),
    .A2(_1746_),
    .B1(_1763_),
    .B2(_1759_),
    .ZN(_1851_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_2 _6622_ (.A1(_1778_),
    .A2(_1845_),
    .B1(_1851_),
    .B2(_1806_),
    .ZN(_1852_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6623_ (.A1(_0671_),
    .A2(_1721_),
    .ZN(_1853_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _6624_ (.I(_1853_),
    .ZN(_1854_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _6625_ (.A1(_1850_),
    .A2(_1852_),
    .A3(_1854_),
    .Z(_1855_));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_1 _6626_ (.A1(_1838_),
    .A2(_1849_),
    .A3(_1855_),
    .ZN(_1856_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _6627_ (.A1(_1837_),
    .A2(_1856_),
    .Z(_1857_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _6628_ (.A1(_1836_),
    .A2(_1857_),
    .ZN(_1858_));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_1 _6629_ (.A1(_1827_),
    .A2(_1833_),
    .A3(_1858_),
    .ZN(_1859_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6630_ (.A1(_1795_),
    .A2(_1859_),
    .ZN(_1860_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _6631_ (.A1(\as2650.r123_2[1][6] ),
    .A2(_1729_),
    .B(_1860_),
    .ZN(_1861_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6632_ (.A1(_1201_),
    .A2(_1717_),
    .ZN(_1862_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6633_ (.A1(_1861_),
    .A2(_1862_),
    .ZN(_0082_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6634_ (.A1(_1833_),
    .A2(_1858_),
    .ZN(_1863_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6635_ (.A1(_1833_),
    .A2(_1858_),
    .ZN(_1864_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _6636_ (.A1(_1827_),
    .A2(_1863_),
    .B(_1864_),
    .ZN(_1865_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _6637_ (.A1(_1837_),
    .A2(_1856_),
    .Z(_1866_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _6638_ (.A1(_1836_),
    .A2(_1857_),
    .B(_1866_),
    .ZN(_1867_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6639_ (.A1(_1852_),
    .A2(_1854_),
    .ZN(_1868_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6640_ (.A1(_1852_),
    .A2(_1854_),
    .ZN(_1869_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6641_ (.A1(_1850_),
    .A2(_1868_),
    .B(_1869_),
    .ZN(_1870_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6642_ (.A1(_1838_),
    .A2(_1849_),
    .ZN(_1871_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6643_ (.A1(_1838_),
    .A2(_1849_),
    .ZN(_1872_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6644_ (.A1(_1871_),
    .A2(_1855_),
    .B(_1872_),
    .ZN(_1873_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6645_ (.A1(_1844_),
    .A2(_1848_),
    .ZN(_1874_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6646_ (.A1(_0671_),
    .A2(_1731_),
    .ZN(_1875_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6647_ (.A1(\as2650.r0[4] ),
    .A2(_1762_),
    .ZN(_1876_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6648_ (.A1(\as2650.r0[5] ),
    .A2(_1745_),
    .ZN(_1877_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _6649_ (.A1(_1876_),
    .A2(_1877_),
    .Z(_1878_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _6650_ (.A1(_1875_),
    .A2(_1878_),
    .Z(_1879_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6651_ (.A1(\as2650.r0[1] ),
    .A2(_1840_),
    .ZN(_1880_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6652_ (.A1(\as2650.r0[2] ),
    .A2(_1809_),
    .ZN(_1881_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _6653_ (.I0(\as2650.r123[0][7] ),
    .I1(\as2650.r123_2[0][7] ),
    .S(_4144_),
    .Z(_1882_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6654_ (.A1(\as2650.r0[0] ),
    .A2(_1882_),
    .ZN(_1883_));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_1 _6655_ (.A1(_1880_),
    .A2(_1881_),
    .A3(_1883_),
    .ZN(_1884_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _6656_ (.A1(_1843_),
    .A2(_1884_),
    .ZN(_1885_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _6657_ (.A1(_1874_),
    .A2(_1879_),
    .A3(_1885_),
    .Z(_1886_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6658_ (.I(_1781_),
    .Z(_1887_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6659_ (.A1(_0364_),
    .A2(_1887_),
    .ZN(_1888_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _6660_ (.A1(_0498_),
    .A2(_1748_),
    .B1(_1783_),
    .B2(_0362_),
    .ZN(_1889_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _6661_ (.A1(_1807_),
    .A2(_1876_),
    .B1(_1889_),
    .B2(_1846_),
    .ZN(_1890_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6662_ (.A1(_4366_),
    .A2(_1720_),
    .ZN(_1891_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _6663_ (.A1(_1890_),
    .A2(_1891_),
    .Z(_1892_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _6664_ (.A1(_1888_),
    .A2(_1892_),
    .ZN(_1893_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _6665_ (.A1(_1886_),
    .A2(_1893_),
    .Z(_1894_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _6666_ (.A1(_1873_),
    .A2(_1894_),
    .Z(_1895_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _6667_ (.A1(_1870_),
    .A2(_1895_),
    .ZN(_1896_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _6668_ (.A1(_1867_),
    .A2(_1896_),
    .ZN(_1897_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _6669_ (.A1(_1865_),
    .A2(_1897_),
    .ZN(_1898_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6670_ (.A1(_1795_),
    .A2(_1898_),
    .ZN(_1899_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _6671_ (.A1(\as2650.r123_2[1][7] ),
    .A2(_1729_),
    .B(_1899_),
    .ZN(_1900_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6672_ (.A1(_1223_),
    .A2(_1717_),
    .ZN(_1901_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6673_ (.A1(_1900_),
    .A2(_1901_),
    .ZN(_0083_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6674_ (.A1(_4467_),
    .A2(_4457_),
    .ZN(_1902_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6675_ (.I(_1902_),
    .Z(_1903_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6676_ (.I(_1903_),
    .Z(_1904_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6677_ (.I(_1904_),
    .Z(_1905_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _6678_ (.A1(_0866_),
    .A2(_1905_),
    .A3(_0960_),
    .ZN(_1906_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6679_ (.I(_1906_),
    .Z(_1907_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6680_ (.I(_1907_),
    .Z(_1908_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6681_ (.I(_1907_),
    .Z(_1909_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6682_ (.A1(\as2650.stack[1][8] ),
    .A2(_1909_),
    .ZN(_1910_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _6683_ (.A1(_1653_),
    .A2(_1908_),
    .B(_1910_),
    .ZN(_0084_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6684_ (.I(_1906_),
    .Z(_1911_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6685_ (.A1(\as2650.stack[1][9] ),
    .A2(_1911_),
    .ZN(_1912_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _6686_ (.A1(_1663_),
    .A2(_1908_),
    .B(_1912_),
    .ZN(_0085_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6687_ (.A1(\as2650.stack[1][10] ),
    .A2(_1911_),
    .ZN(_1913_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _6688_ (.A1(_1666_),
    .A2(_1908_),
    .B(_1913_),
    .ZN(_0086_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6689_ (.A1(\as2650.stack[1][11] ),
    .A2(_1911_),
    .ZN(_1914_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _6690_ (.A1(_1668_),
    .A2(_1908_),
    .B(_1914_),
    .ZN(_0087_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6691_ (.A1(\as2650.stack[1][12] ),
    .A2(_1911_),
    .ZN(_1915_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _6692_ (.A1(_1670_),
    .A2(_1909_),
    .B(_1915_),
    .ZN(_0088_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6693_ (.A1(\as2650.stack[1][13] ),
    .A2(_1907_),
    .ZN(_1916_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _6694_ (.A1(_1672_),
    .A2(_1909_),
    .B(_1916_),
    .ZN(_0089_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6695_ (.A1(\as2650.stack[1][14] ),
    .A2(_1907_),
    .ZN(_1917_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _6696_ (.A1(_1674_),
    .A2(_1909_),
    .B(_1917_),
    .ZN(_0090_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6697_ (.A1(_4456_),
    .A2(_4458_),
    .ZN(_1918_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6698_ (.I(_1918_),
    .Z(_1919_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6699_ (.I(_1919_),
    .Z(_1920_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6700_ (.I(_1920_),
    .Z(_1921_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _6701_ (.A1(_0866_),
    .A2(_1921_),
    .A3(_0960_),
    .ZN(_1922_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6702_ (.I(_1922_),
    .Z(_1923_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6703_ (.I(_1923_),
    .Z(_1924_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6704_ (.I(_1923_),
    .Z(_1925_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6705_ (.A1(\as2650.stack[0][8] ),
    .A2(_1925_),
    .ZN(_1926_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _6706_ (.A1(_1653_),
    .A2(_1924_),
    .B(_1926_),
    .ZN(_0091_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6707_ (.I(_1922_),
    .Z(_1927_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6708_ (.A1(\as2650.stack[0][9] ),
    .A2(_1927_),
    .ZN(_1928_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _6709_ (.A1(_1663_),
    .A2(_1924_),
    .B(_1928_),
    .ZN(_0092_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6710_ (.A1(\as2650.stack[0][10] ),
    .A2(_1927_),
    .ZN(_1929_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _6711_ (.A1(_1666_),
    .A2(_1924_),
    .B(_1929_),
    .ZN(_0093_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6712_ (.A1(\as2650.stack[0][11] ),
    .A2(_1927_),
    .ZN(_1930_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _6713_ (.A1(_1668_),
    .A2(_1924_),
    .B(_1930_),
    .ZN(_0094_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6714_ (.A1(\as2650.stack[0][12] ),
    .A2(_1927_),
    .ZN(_1931_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _6715_ (.A1(_1670_),
    .A2(_1925_),
    .B(_1931_),
    .ZN(_0095_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6716_ (.A1(\as2650.stack[0][13] ),
    .A2(_1923_),
    .ZN(_1932_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _6717_ (.A1(_1672_),
    .A2(_1925_),
    .B(_1932_),
    .ZN(_0096_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6718_ (.A1(\as2650.stack[0][14] ),
    .A2(_1923_),
    .ZN(_1933_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _6719_ (.A1(_1674_),
    .A2(_1925_),
    .B(_1933_),
    .ZN(_0097_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _6720_ (.A1(_1059_),
    .A2(_1145_),
    .A3(_1165_),
    .ZN(_1934_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6721_ (.A1(_4195_),
    .A2(_1164_),
    .ZN(_1935_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _6722_ (.A1(_1038_),
    .A2(_1215_),
    .A3(_1133_),
    .A4(_1935_),
    .ZN(_1936_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6723_ (.A1(_1934_),
    .A2(_1936_),
    .B(_1261_),
    .ZN(_1937_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6724_ (.I(_1937_),
    .Z(_1938_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _6725_ (.I(_1716_),
    .Z(_1939_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6726_ (.A1(_1612_),
    .A2(_1051_),
    .ZN(_1940_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _6727_ (.A1(_1939_),
    .A2(_1035_),
    .B(_1940_),
    .C(_4438_),
    .ZN(_1941_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6728_ (.I(_1941_),
    .Z(_1942_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _6729_ (.A1(_1867_),
    .A2(_1896_),
    .Z(_1943_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6730_ (.A1(_1865_),
    .A2(_1897_),
    .B(_1943_),
    .ZN(_1944_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6731_ (.A1(_1873_),
    .A2(_1894_),
    .ZN(_1945_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6732_ (.A1(_1870_),
    .A2(_1895_),
    .ZN(_1946_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6733_ (.A1(_1945_),
    .A2(_1946_),
    .ZN(_1947_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _6734_ (.A1(_0788_),
    .A2(_1736_),
    .A3(_1890_),
    .ZN(_1948_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6735_ (.A1(_1888_),
    .A2(_1892_),
    .B(_1948_),
    .ZN(_1949_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6736_ (.A1(_1879_),
    .A2(_1885_),
    .ZN(_1950_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _6737_ (.A1(_1879_),
    .A2(_1885_),
    .Z(_1951_));
 gf180mcu_fd_sc_mcu7t5v0__oai32_1 _6738_ (.A1(_1874_),
    .A2(_1950_),
    .A3(_1951_),
    .B1(_1886_),
    .B2(_1893_),
    .ZN(_1952_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6739_ (.A1(\as2650.r0[5] ),
    .A2(_1761_),
    .ZN(_1953_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _6740_ (.A1(_1847_),
    .A2(_1953_),
    .Z(_1954_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _6741_ (.A1(_0672_),
    .A2(_1732_),
    .A3(_1878_),
    .ZN(_1955_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _6742_ (.A1(_1954_),
    .A2(_1955_),
    .Z(_1956_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6743_ (.A1(_0499_),
    .A2(_1887_),
    .ZN(_1957_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _6744_ (.A1(_1956_),
    .A2(_1957_),
    .ZN(_1958_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6745_ (.A1(_1843_),
    .A2(_1884_),
    .ZN(_1959_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6746_ (.A1(_1879_),
    .A2(_1885_),
    .B(_1959_),
    .ZN(_1960_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6747_ (.A1(\as2650.r0[7] ),
    .A2(_1730_),
    .ZN(_1961_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6748_ (.A1(\as2650.r0[6] ),
    .A2(_1744_),
    .ZN(_1962_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _6749_ (.A1(_1953_),
    .A2(_1962_),
    .ZN(_1963_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _6750_ (.A1(_1961_),
    .A2(_1963_),
    .ZN(_1964_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6751_ (.I(_1882_),
    .Z(_1965_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6752_ (.A1(\as2650.r0[1] ),
    .A2(_1965_),
    .ZN(_1966_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _6753_ (.A1(_1880_),
    .A2(_1883_),
    .Z(_1967_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_2 _6754_ (.A1(_1842_),
    .A2(_1966_),
    .B1(_1967_),
    .B2(_1881_),
    .ZN(_1968_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6755_ (.A1(\as2650.r0[3] ),
    .A2(_1810_),
    .ZN(_1969_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6756_ (.I(_1840_),
    .Z(_1970_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6757_ (.A1(_4519_),
    .A2(_1970_),
    .ZN(_1971_));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_1 _6758_ (.A1(_1966_),
    .A2(_1969_),
    .A3(_1971_),
    .ZN(_1972_));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_1 _6759_ (.A1(_1964_),
    .A2(_1968_),
    .A3(_1972_),
    .ZN(_1973_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _6760_ (.A1(_1960_),
    .A2(_1973_),
    .ZN(_1974_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _6761_ (.A1(_1958_),
    .A2(_1974_),
    .Z(_1975_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _6762_ (.A1(_1952_),
    .A2(_1975_),
    .Z(_1976_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _6763_ (.A1(_1949_),
    .A2(_1976_),
    .ZN(_1977_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _6764_ (.A1(_1947_),
    .A2(_1977_),
    .ZN(_1978_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _6765_ (.A1(_1944_),
    .A2(_1978_),
    .Z(_1979_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6766_ (.I(_1741_),
    .Z(_1980_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _6767_ (.A1(\as2650.r123_2[2][0] ),
    .A2(_1942_),
    .B1(_1979_),
    .B2(_1980_),
    .ZN(_1981_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6768_ (.A1(_1713_),
    .A2(_1938_),
    .B(_1981_),
    .ZN(_0098_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _6769_ (.A1(_1116_),
    .A2(_1940_),
    .B1(_1942_),
    .B2(\as2650.r123_2[2][1] ),
    .ZN(_1982_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _6770_ (.A1(_1945_),
    .A2(_1946_),
    .B(_1977_),
    .ZN(_1983_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _6771_ (.A1(_1944_),
    .A2(_1978_),
    .B(_1983_),
    .ZN(_1984_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _6772_ (.A1(_1952_),
    .A2(_1975_),
    .Z(_1985_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _6773_ (.A1(_1949_),
    .A2(_1976_),
    .B(_1985_),
    .ZN(_1986_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _6774_ (.A1(_1956_),
    .A2(_1957_),
    .Z(_1987_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6775_ (.A1(_1960_),
    .A2(_1973_),
    .ZN(_1988_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6776_ (.A1(_1958_),
    .A2(_1974_),
    .B(_1988_),
    .ZN(_1989_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6777_ (.A1(_1953_),
    .A2(_1962_),
    .ZN(_1990_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6778_ (.A1(_1961_),
    .A2(_1963_),
    .ZN(_1991_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6779_ (.A1(_1990_),
    .A2(_1991_),
    .ZN(_1992_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6780_ (.A1(_0586_),
    .A2(_1887_),
    .ZN(_1993_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _6781_ (.A1(_1992_),
    .A2(_1993_),
    .Z(_1994_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6782_ (.A1(_1992_),
    .A2(_1993_),
    .ZN(_1995_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6783_ (.A1(_1994_),
    .A2(_1995_),
    .ZN(_1996_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6784_ (.A1(_1968_),
    .A2(_1972_),
    .ZN(_1997_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6785_ (.A1(_1968_),
    .A2(_1972_),
    .ZN(_1998_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6786_ (.A1(_1964_),
    .A2(_1997_),
    .B(_1998_),
    .ZN(_1999_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _6787_ (.A1(_4366_),
    .A2(_1749_),
    .B1(_1764_),
    .B2(_0672_),
    .ZN(_2000_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6788_ (.A1(_4366_),
    .A2(_1763_),
    .ZN(_2001_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6789_ (.A1(_1962_),
    .A2(_2001_),
    .ZN(_2002_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6790_ (.A1(_2000_),
    .A2(_2002_),
    .ZN(_2003_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6791_ (.A1(_4519_),
    .A2(_1965_),
    .ZN(_2004_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6792_ (.I(_1965_),
    .Z(_2005_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _6793_ (.A1(_1757_),
    .A2(_2005_),
    .B1(_1970_),
    .B2(_4520_),
    .ZN(_2006_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _6794_ (.A1(_1880_),
    .A2(_2004_),
    .B1(_2006_),
    .B2(_1969_),
    .ZN(_2007_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6795_ (.A1(_0362_),
    .A2(_1841_),
    .ZN(_2008_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _6796_ (.A1(_0498_),
    .A2(_1811_),
    .Z(_2009_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _6797_ (.A1(_2004_),
    .A2(_2008_),
    .A3(_2009_),
    .Z(_2010_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _6798_ (.A1(_2007_),
    .A2(_2010_),
    .Z(_2011_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _6799_ (.A1(_2003_),
    .A2(_2011_),
    .Z(_2012_));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_1 _6800_ (.A1(_1996_),
    .A2(_1999_),
    .A3(_2012_),
    .ZN(_2013_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _6801_ (.A1(_1989_),
    .A2(_2013_),
    .ZN(_2014_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _6802_ (.A1(_1987_),
    .A2(_2014_),
    .ZN(_2015_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _6803_ (.A1(_1986_),
    .A2(_2015_),
    .ZN(_2016_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _6804_ (.A1(_1984_),
    .A2(_2016_),
    .Z(_2017_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6805_ (.A1(_1727_),
    .A2(_2017_),
    .ZN(_2018_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6806_ (.A1(_1982_),
    .A2(_2018_),
    .ZN(_0099_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6807_ (.I(_1941_),
    .Z(_2019_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _6808_ (.A1(_1986_),
    .A2(_2015_),
    .Z(_2020_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _6809_ (.A1(_1984_),
    .A2(_2016_),
    .B(_2020_),
    .ZN(_2021_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6810_ (.A1(_1989_),
    .A2(_2013_),
    .ZN(_2022_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6811_ (.A1(_1987_),
    .A2(_2014_),
    .B(_2022_),
    .ZN(_2023_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6812_ (.A1(_1999_),
    .A2(_2012_),
    .ZN(_2024_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6813_ (.A1(_1999_),
    .A2(_2012_),
    .ZN(_2025_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6814_ (.A1(_1996_),
    .A2(_2024_),
    .B(_2025_),
    .ZN(_2026_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6815_ (.I(_1887_),
    .Z(_2027_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _6816_ (.A1(_2027_),
    .A2(_2002_),
    .Z(_2028_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _6817_ (.A1(_0750_),
    .A2(_2027_),
    .B(_2002_),
    .ZN(_2029_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6818_ (.A1(_2028_),
    .A2(_2029_),
    .ZN(_2030_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6819_ (.A1(_2007_),
    .A2(_2010_),
    .ZN(_2031_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6820_ (.A1(_2003_),
    .A2(_2011_),
    .ZN(_2032_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6821_ (.A1(_2031_),
    .A2(_2032_),
    .ZN(_2033_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6822_ (.A1(_2004_),
    .A2(_2008_),
    .ZN(_2034_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6823_ (.A1(_0362_),
    .A2(_1965_),
    .ZN(_2035_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6824_ (.A1(_1971_),
    .A2(_2035_),
    .ZN(_2036_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _6825_ (.A1(_2034_),
    .A2(_2009_),
    .B(_2036_),
    .ZN(_2037_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6826_ (.A1(\as2650.r0[4] ),
    .A2(_1841_),
    .ZN(_2038_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _6827_ (.A1(_0585_),
    .A2(_1810_),
    .Z(_2039_));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_1 _6828_ (.A1(_2035_),
    .A2(_2038_),
    .A3(_2039_),
    .ZN(_2040_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _6829_ (.A1(_2037_),
    .A2(_2040_),
    .Z(_2041_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _6830_ (.A1(_2001_),
    .A2(_2041_),
    .Z(_2042_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _6831_ (.A1(_2033_),
    .A2(_2042_),
    .ZN(_2043_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _6832_ (.A1(_2030_),
    .A2(_2043_),
    .Z(_2044_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _6833_ (.A1(_2026_),
    .A2(_2044_),
    .ZN(_2045_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _6834_ (.A1(_1994_),
    .A2(_2045_),
    .Z(_2046_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _6835_ (.A1(_2023_),
    .A2(_2046_),
    .Z(_2047_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _6836_ (.A1(_2021_),
    .A2(_2047_),
    .Z(_2048_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _6837_ (.A1(\as2650.r123_2[2][2] ),
    .A2(_2019_),
    .B1(_2048_),
    .B2(_1980_),
    .ZN(_2049_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6838_ (.A1(_1139_),
    .A2(_1938_),
    .B(_2049_),
    .ZN(_0100_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _6839_ (.A1(_2023_),
    .A2(_2046_),
    .Z(_2050_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _6840_ (.A1(_2021_),
    .A2(_2047_),
    .B(_2050_),
    .ZN(_2051_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6841_ (.A1(_2026_),
    .A2(_2044_),
    .ZN(_2052_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _6842_ (.A1(_1994_),
    .A2(_2045_),
    .Z(_2053_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _6843_ (.I(_2042_),
    .ZN(_2054_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6844_ (.A1(_2033_),
    .A2(_2054_),
    .ZN(_2055_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6845_ (.A1(_2030_),
    .A2(_2043_),
    .ZN(_2056_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6846_ (.A1(_2055_),
    .A2(_2056_),
    .ZN(_2057_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6847_ (.A1(_0788_),
    .A2(_2027_),
    .ZN(_2058_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6848_ (.A1(_0499_),
    .A2(_2005_),
    .ZN(_2059_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _6849_ (.A1(_0671_),
    .A2(_1811_),
    .Z(_2060_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6850_ (.A1(_0585_),
    .A2(_1970_),
    .ZN(_2061_));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_1 _6851_ (.A1(_2059_),
    .A2(_2060_),
    .A3(_2061_),
    .ZN(_2062_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6852_ (.A1(_2035_),
    .A2(_2038_),
    .ZN(_2063_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6853_ (.A1(_2008_),
    .A2(_2059_),
    .ZN(_2064_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _6854_ (.A1(_2063_),
    .A2(_2039_),
    .B(_2064_),
    .ZN(_2065_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _6855_ (.A1(_2062_),
    .A2(_2065_),
    .Z(_2066_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _6856_ (.A1(_4367_),
    .A2(_1764_),
    .A3(_2041_),
    .ZN(_2067_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6857_ (.A1(_2037_),
    .A2(_2040_),
    .B(_2067_),
    .ZN(_2068_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _6858_ (.A1(_2066_),
    .A2(_2068_),
    .ZN(_2069_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _6859_ (.A1(_2058_),
    .A2(_2069_),
    .Z(_2070_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _6860_ (.A1(_2057_),
    .A2(_2070_),
    .Z(_2071_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _6861_ (.A1(_2028_),
    .A2(_2071_),
    .ZN(_2072_));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _6862_ (.A1(_2052_),
    .A2(_2053_),
    .A3(_2072_),
    .Z(_2073_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _6863_ (.A1(_2052_),
    .A2(_2053_),
    .B(_2072_),
    .ZN(_2074_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6864_ (.A1(_2073_),
    .A2(_2074_),
    .ZN(_2075_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _6865_ (.A1(_2051_),
    .A2(_2075_),
    .ZN(_2076_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _6866_ (.A1(\as2650.r123_2[2][3] ),
    .A2(_2019_),
    .B1(_2076_),
    .B2(_1980_),
    .ZN(_2077_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6867_ (.A1(_1156_),
    .A2(_1938_),
    .B(_2077_),
    .ZN(_0101_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _6868_ (.A1(_2062_),
    .A2(_2065_),
    .Z(_2078_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _6869_ (.I(_2078_),
    .ZN(_2079_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6870_ (.A1(_2059_),
    .A2(_2061_),
    .ZN(_2080_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6871_ (.A1(_2059_),
    .A2(_2061_),
    .ZN(_2081_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _6872_ (.A1(_2060_),
    .A2(_2080_),
    .B(_2081_),
    .ZN(_2082_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6873_ (.A1(_0586_),
    .A2(_2005_),
    .ZN(_2083_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _6874_ (.I(_1970_),
    .Z(_2084_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6875_ (.A1(_0750_),
    .A2(_2084_),
    .ZN(_2085_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _6876_ (.A1(_2083_),
    .A2(_2085_),
    .ZN(_2086_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6877_ (.A1(_4367_),
    .A2(_1812_),
    .ZN(_2087_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _6878_ (.A1(_2086_),
    .A2(_2087_),
    .ZN(_2088_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _6879_ (.A1(_2082_),
    .A2(_2088_),
    .Z(_2089_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _6880_ (.A1(_2079_),
    .A2(_2089_),
    .Z(_2090_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6881_ (.A1(_2066_),
    .A2(_2068_),
    .ZN(_2091_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6882_ (.A1(_2058_),
    .A2(_2069_),
    .B(_2091_),
    .ZN(_2092_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _6883_ (.A1(_2090_),
    .A2(_2092_),
    .Z(_2093_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6884_ (.A1(_2057_),
    .A2(_2070_),
    .ZN(_2094_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6885_ (.A1(_2028_),
    .A2(_2071_),
    .ZN(_2095_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6886_ (.A1(_2094_),
    .A2(_2095_),
    .ZN(_2096_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _6887_ (.A1(_2093_),
    .A2(_2096_),
    .ZN(_2097_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_2 _6888_ (.A1(_2021_),
    .A2(_2047_),
    .B(_2074_),
    .C(_2050_),
    .ZN(_2098_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6889_ (.A1(_2073_),
    .A2(_2098_),
    .ZN(_2099_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _6890_ (.A1(_2097_),
    .A2(_2099_),
    .Z(_2100_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6891_ (.A1(_1794_),
    .A2(_2100_),
    .ZN(_2101_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _6892_ (.A1(\as2650.r123_2[2][4] ),
    .A2(_1942_),
    .B(_2101_),
    .ZN(_2102_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6893_ (.A1(_1174_),
    .A2(_1938_),
    .B(_2102_),
    .ZN(_0102_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6894_ (.A1(_2090_),
    .A2(_2092_),
    .ZN(_2103_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6895_ (.A1(_2093_),
    .A2(_2096_),
    .ZN(_2104_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_1 _6896_ (.A1(_2073_),
    .A2(_2097_),
    .A3(_2098_),
    .B(_2104_),
    .ZN(_2105_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _6897_ (.A1(_2082_),
    .A2(_2088_),
    .Z(_2106_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6898_ (.A1(_2079_),
    .A2(_2089_),
    .ZN(_2107_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6899_ (.A1(_2106_),
    .A2(_2107_),
    .ZN(_2108_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6900_ (.I(_2005_),
    .Z(_2109_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6901_ (.A1(_0750_),
    .A2(_2109_),
    .ZN(_2110_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _6902_ (.A1(_2061_),
    .A2(_2110_),
    .B1(_2086_),
    .B2(_2087_),
    .ZN(_2111_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6903_ (.A1(_0788_),
    .A2(_2084_),
    .ZN(_2112_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _6904_ (.A1(_2110_),
    .A2(_2112_),
    .Z(_2113_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _6905_ (.A1(_2111_),
    .A2(_2113_),
    .ZN(_2114_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _6906_ (.A1(_2108_),
    .A2(_2114_),
    .ZN(_2115_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _6907_ (.I(_2115_),
    .ZN(_2116_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _6908_ (.A1(_2103_),
    .A2(_2105_),
    .A3(_2116_),
    .Z(_2117_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _6909_ (.A1(\as2650.r123_2[2][5] ),
    .A2(_2019_),
    .B1(_2117_),
    .B2(_1980_),
    .ZN(_2118_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6910_ (.A1(_1189_),
    .A2(_1937_),
    .B(_2118_),
    .ZN(_0103_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _6911_ (.A1(_1201_),
    .A2(_1940_),
    .B1(_1942_),
    .B2(\as2650.r123_2[2][6] ),
    .ZN(_2119_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6912_ (.A1(_2103_),
    .A2(_2116_),
    .ZN(_2120_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6913_ (.A1(_2103_),
    .A2(_2116_),
    .ZN(_2121_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _6914_ (.A1(_2105_),
    .A2(_2120_),
    .B(_2121_),
    .ZN(_2122_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6915_ (.A1(_2107_),
    .A2(_2114_),
    .ZN(_2123_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _6916_ (.A1(_0789_),
    .A2(_2109_),
    .A3(_2085_),
    .ZN(_2124_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6917_ (.A1(_2111_),
    .A2(_2113_),
    .ZN(_2125_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6918_ (.A1(_2106_),
    .A2(_2114_),
    .B(_2125_),
    .ZN(_2126_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _6919_ (.A1(_2124_),
    .A2(_2126_),
    .Z(_2127_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _6920_ (.A1(_2123_),
    .A2(_2127_),
    .Z(_2128_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _6921_ (.A1(_2122_),
    .A2(_2128_),
    .Z(_2129_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6922_ (.A1(_1727_),
    .A2(_2129_),
    .ZN(_2130_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6923_ (.A1(_2119_),
    .A2(_2130_),
    .ZN(_0104_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _6924_ (.A1(_2107_),
    .A2(_2114_),
    .A3(_2127_),
    .ZN(_2131_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6925_ (.A1(_2122_),
    .A2(_2128_),
    .ZN(_2132_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6926_ (.A1(_0791_),
    .A2(_2109_),
    .ZN(_2133_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _6927_ (.A1(_0752_),
    .A2(_2084_),
    .B(_2126_),
    .ZN(_2134_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6928_ (.A1(_2133_),
    .A2(_2134_),
    .ZN(_2135_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _6929_ (.A1(_2131_),
    .A2(_2132_),
    .A3(_2135_),
    .ZN(_2136_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _6930_ (.A1(_1223_),
    .A2(_1940_),
    .B1(_2019_),
    .B2(\as2650.r123_2[2][7] ),
    .ZN(_2137_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6931_ (.A1(_1795_),
    .A2(_2136_),
    .B(_2137_),
    .ZN(_0105_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6932_ (.I(_4295_),
    .Z(_2138_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6933_ (.I(_0850_),
    .Z(_2139_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6934_ (.A1(_2139_),
    .A2(_1640_),
    .ZN(_2140_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _6935_ (.A1(_0967_),
    .A2(_2140_),
    .Z(_2141_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6936_ (.I(_2141_),
    .Z(_2142_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6937_ (.I(_2142_),
    .Z(_2143_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6938_ (.I(_0862_),
    .Z(_2144_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _6939_ (.I(_2144_),
    .Z(_2145_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6940_ (.I(_2145_),
    .Z(_2146_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6941_ (.I(_2146_),
    .Z(_2147_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6942_ (.I(_0957_),
    .Z(_2148_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6943_ (.I(_0873_),
    .Z(_2149_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _6944_ (.I(_0868_),
    .Z(_2150_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6945_ (.A1(_2150_),
    .A2(_4176_),
    .ZN(_2151_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6946_ (.A1(_1335_),
    .A2(_2151_),
    .ZN(_2152_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _6947_ (.I(_0881_),
    .Z(_2153_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6948_ (.I(_0895_),
    .Z(_2154_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _6949_ (.A1(_1500_),
    .A2(_1309_),
    .B(_2154_),
    .ZN(_2155_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6950_ (.A1(_0868_),
    .A2(_1682_),
    .ZN(_2156_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _6951_ (.I(_2156_),
    .Z(_2157_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _6952_ (.A1(_2153_),
    .A2(_0889_),
    .B(_2155_),
    .C(_2157_),
    .ZN(_2158_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6953_ (.A1(_2152_),
    .A2(_2158_),
    .ZN(_2159_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6954_ (.I(_0898_),
    .Z(_2160_));
 gf180mcu_fd_sc_mcu7t5v0__oai32_1 _6955_ (.A1(_2149_),
    .A2(_0875_),
    .A3(_2159_),
    .B1(_0897_),
    .B2(_2160_),
    .ZN(_2161_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6956_ (.A1(_0969_),
    .A2(_2161_),
    .ZN(_2162_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _6957_ (.A1(_2148_),
    .A2(_1657_),
    .A3(_2162_),
    .ZN(_2163_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6958_ (.I(_2163_),
    .Z(_2164_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6959_ (.I(_0900_),
    .Z(_2165_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6960_ (.A1(_2139_),
    .A2(_1657_),
    .ZN(_2166_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6961_ (.A1(_2165_),
    .A2(_2166_),
    .ZN(_2167_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6962_ (.I(_2167_),
    .Z(_2168_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _6963_ (.A1(_2147_),
    .A2(_2164_),
    .B1(_2168_),
    .B2(\as2650.stack[2][0] ),
    .C(_2142_),
    .ZN(_2169_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _6964_ (.A1(_2138_),
    .A2(_2143_),
    .B(_2169_),
    .ZN(_0106_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _6965_ (.I(_0912_),
    .Z(_2170_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6966_ (.I(_2163_),
    .Z(_2171_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6967_ (.I(_2167_),
    .Z(_2172_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6968_ (.I(_2141_),
    .Z(_2173_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _6969_ (.A1(_2170_),
    .A2(_2171_),
    .B1(_2172_),
    .B2(\as2650.stack[2][1] ),
    .C(_2173_),
    .ZN(_2174_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6970_ (.I(_0858_),
    .Z(_2175_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6971_ (.A1(_2175_),
    .A2(_2140_),
    .ZN(_2176_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6972_ (.A1(_0908_),
    .A2(_2176_),
    .ZN(_2177_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6973_ (.A1(_2174_),
    .A2(_2177_),
    .ZN(_0107_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _6974_ (.I(_0920_),
    .Z(_2178_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _6975_ (.A1(_2178_),
    .A2(_2171_),
    .B1(_2172_),
    .B2(\as2650.stack[2][2] ),
    .C(_2173_),
    .ZN(_2179_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6976_ (.A1(_0918_),
    .A2(_2176_),
    .ZN(_2180_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6977_ (.A1(_2179_),
    .A2(_2180_),
    .ZN(_0108_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _6978_ (.I(\as2650.pc[3] ),
    .Z(_2181_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6979_ (.I(_2181_),
    .Z(_2182_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _6980_ (.I(_2182_),
    .Z(_2183_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _6981_ (.A1(_2183_),
    .A2(_2171_),
    .B1(_2172_),
    .B2(\as2650.stack[2][3] ),
    .C(_2173_),
    .ZN(_2184_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6982_ (.A1(_0925_),
    .A2(_2176_),
    .ZN(_2185_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6983_ (.A1(_2184_),
    .A2(_2185_),
    .ZN(_0109_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6984_ (.I(_0617_),
    .Z(_2186_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _6985_ (.I(\as2650.pc[4] ),
    .Z(_2187_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _6986_ (.I(_2187_),
    .Z(_2188_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6987_ (.I(_2188_),
    .Z(_2189_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _6988_ (.I(_2189_),
    .Z(_2190_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _6989_ (.I(_2190_),
    .Z(_2191_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _6990_ (.A1(_2191_),
    .A2(_2164_),
    .B1(_2168_),
    .B2(\as2650.stack[2][4] ),
    .C(_2142_),
    .ZN(_2192_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _6991_ (.A1(_2186_),
    .A2(_2143_),
    .B(_2192_),
    .ZN(_0110_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6992_ (.I(_0937_),
    .Z(_2193_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _6993_ (.I(\as2650.pc[5] ),
    .Z(_2194_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6994_ (.I(_2194_),
    .Z(_2195_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6995_ (.I(_2195_),
    .Z(_2196_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _6996_ (.I(_2196_),
    .Z(_2197_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _6997_ (.A1(_2197_),
    .A2(_2164_),
    .B1(_2168_),
    .B2(\as2650.stack[2][5] ),
    .C(_2142_),
    .ZN(_2198_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _6998_ (.A1(_2193_),
    .A2(_2143_),
    .B(_2198_),
    .ZN(_0111_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6999_ (.I(_1530_),
    .Z(_2199_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7000_ (.I(_2199_),
    .Z(_2200_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _7001_ (.I(_0947_),
    .Z(_2201_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _7002_ (.A1(_2201_),
    .A2(_2164_),
    .B1(_2168_),
    .B2(\as2650.stack[2][6] ),
    .C(_2173_),
    .ZN(_2202_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _7003_ (.A1(_2200_),
    .A2(_2143_),
    .B(_2202_),
    .ZN(_0112_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _7004_ (.I(\as2650.pc[7] ),
    .Z(_2203_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7005_ (.I(_2203_),
    .Z(_2204_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _7006_ (.I(_2204_),
    .Z(_2205_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _7007_ (.A1(_2205_),
    .A2(_2171_),
    .B1(_2172_),
    .B2(\as2650.stack[2][7] ),
    .C(_2141_),
    .ZN(_2206_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _7008_ (.A1(_0951_),
    .A2(_2176_),
    .ZN(_2207_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _7009_ (.A1(_2206_),
    .A2(_2207_),
    .ZN(_0113_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7010_ (.A1(_1118_),
    .A2(_1009_),
    .ZN(_2208_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _7011_ (.A1(_1018_),
    .A2(_2208_),
    .ZN(_2209_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7012_ (.I(_2209_),
    .Z(_2210_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7013_ (.I(_2210_),
    .Z(_2211_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7014_ (.I(_2162_),
    .Z(_2212_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _7015_ (.A1(_0622_),
    .A2(_2212_),
    .ZN(_2213_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7016_ (.I(_2213_),
    .Z(_2214_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7017_ (.I(_4474_),
    .Z(_2215_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7018_ (.A1(_2215_),
    .A2(_0901_),
    .ZN(_2216_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7019_ (.I(_2216_),
    .Z(_2217_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _7020_ (.A1(_2147_),
    .A2(_2214_),
    .B1(_2217_),
    .B2(\as2650.stack[4][0] ),
    .C(_2210_),
    .ZN(_2218_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _7021_ (.A1(_2138_),
    .A2(_2211_),
    .B(_2218_),
    .ZN(_0114_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7022_ (.I(_2213_),
    .Z(_2219_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7023_ (.I(_2216_),
    .Z(_2220_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7024_ (.I(_2209_),
    .Z(_2221_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _7025_ (.A1(_2170_),
    .A2(_2219_),
    .B1(_2220_),
    .B2(\as2650.stack[4][1] ),
    .C(_2221_),
    .ZN(_2222_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _7026_ (.I(_0957_),
    .Z(_2223_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _7027_ (.A1(_2223_),
    .A2(_4482_),
    .A3(_0968_),
    .ZN(_2224_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _7028_ (.A1(_0908_),
    .A2(_2224_),
    .ZN(_2225_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _7029_ (.A1(_2222_),
    .A2(_2225_),
    .ZN(_0115_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _7030_ (.A1(_2178_),
    .A2(_2219_),
    .B1(_2220_),
    .B2(\as2650.stack[4][2] ),
    .C(_2221_),
    .ZN(_2226_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _7031_ (.A1(_0918_),
    .A2(_2224_),
    .ZN(_2227_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _7032_ (.A1(_2226_),
    .A2(_2227_),
    .ZN(_0116_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _7033_ (.A1(_2183_),
    .A2(_2219_),
    .B1(_2220_),
    .B2(\as2650.stack[4][3] ),
    .C(_2221_),
    .ZN(_2228_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _7034_ (.A1(_0925_),
    .A2(_2224_),
    .ZN(_2229_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _7035_ (.A1(_2228_),
    .A2(_2229_),
    .ZN(_0117_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _7036_ (.A1(_2191_),
    .A2(_2214_),
    .B1(_2217_),
    .B2(\as2650.stack[4][4] ),
    .C(_2210_),
    .ZN(_2230_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _7037_ (.A1(_2186_),
    .A2(_2211_),
    .B(_2230_),
    .ZN(_0118_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _7038_ (.A1(_2197_),
    .A2(_2214_),
    .B1(_2217_),
    .B2(\as2650.stack[4][5] ),
    .C(_2210_),
    .ZN(_2231_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _7039_ (.A1(_2193_),
    .A2(_2211_),
    .B(_2231_),
    .ZN(_0119_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _7040_ (.A1(_2201_),
    .A2(_2214_),
    .B1(_2217_),
    .B2(\as2650.stack[4][6] ),
    .C(_2221_),
    .ZN(_2232_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _7041_ (.A1(_2200_),
    .A2(_2211_),
    .B(_2232_),
    .ZN(_0120_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _7042_ (.A1(_2205_),
    .A2(_2219_),
    .B1(_2220_),
    .B2(\as2650.stack[4][7] ),
    .C(_2209_),
    .ZN(_2233_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _7043_ (.A1(_0951_),
    .A2(_2224_),
    .ZN(_2234_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _7044_ (.A1(_2233_),
    .A2(_2234_),
    .ZN(_0121_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7045_ (.I(\as2650.r123_2[3][0] ),
    .Z(_2235_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7046_ (.I(_2235_),
    .Z(_0122_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7047_ (.I(\as2650.r123_2[3][1] ),
    .Z(_2236_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7048_ (.I(_2236_),
    .Z(_0123_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7049_ (.I(\as2650.r123_2[3][2] ),
    .Z(_2237_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7050_ (.I(_2237_),
    .Z(_0124_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7051_ (.I(\as2650.r123_2[3][3] ),
    .Z(_2238_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7052_ (.I(_2238_),
    .Z(_0125_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7053_ (.I(\as2650.r123_2[3][4] ),
    .Z(_2239_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7054_ (.I(_2239_),
    .Z(_0126_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7055_ (.I(\as2650.r123_2[3][5] ),
    .Z(_2240_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7056_ (.I(_2240_),
    .Z(_0127_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7057_ (.I(\as2650.r123_2[3][6] ),
    .Z(_2241_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7058_ (.I(_2241_),
    .Z(_0128_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7059_ (.I(\as2650.r123_2[3][7] ),
    .Z(_2242_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7060_ (.I(_2242_),
    .Z(_0129_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _7061_ (.A1(_0967_),
    .A2(_2166_),
    .Z(_2243_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7062_ (.I(_2243_),
    .Z(_2244_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7063_ (.I(_2244_),
    .Z(_2245_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _7064_ (.A1(_2148_),
    .A2(_1905_),
    .A3(_2162_),
    .ZN(_2246_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7065_ (.I(_2246_),
    .Z(_2247_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _7066_ (.A1(_2139_),
    .A2(_1905_),
    .ZN(_2248_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7067_ (.A1(_2165_),
    .A2(_2248_),
    .ZN(_2249_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7068_ (.I(_2249_),
    .Z(_2250_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _7069_ (.A1(_2147_),
    .A2(_2247_),
    .B1(_2250_),
    .B2(\as2650.stack[1][0] ),
    .C(_2244_),
    .ZN(_2251_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _7070_ (.A1(_2138_),
    .A2(_2245_),
    .B(_2251_),
    .ZN(_0130_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7071_ (.I(_2246_),
    .Z(_2252_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7072_ (.I(_2249_),
    .Z(_2253_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7073_ (.I(_2243_),
    .Z(_2254_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _7074_ (.A1(_2170_),
    .A2(_2252_),
    .B1(_2253_),
    .B2(\as2650.stack[1][1] ),
    .C(_2254_),
    .ZN(_2255_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7075_ (.A1(_2175_),
    .A2(_2166_),
    .ZN(_2256_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _7076_ (.A1(_0908_),
    .A2(_2256_),
    .ZN(_2257_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _7077_ (.A1(_2255_),
    .A2(_2257_),
    .ZN(_0131_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7078_ (.I(_0921_),
    .Z(_2258_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _7079_ (.A1(_2258_),
    .A2(_2252_),
    .B1(_2253_),
    .B2(\as2650.stack[1][2] ),
    .C(_2254_),
    .ZN(_2259_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _7080_ (.A1(_0918_),
    .A2(_2256_),
    .ZN(_2260_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _7081_ (.A1(_2259_),
    .A2(_2260_),
    .ZN(_0132_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _7082_ (.A1(_2183_),
    .A2(_2252_),
    .B1(_2253_),
    .B2(\as2650.stack[1][3] ),
    .C(_2254_),
    .ZN(_2261_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _7083_ (.A1(_0925_),
    .A2(_2256_),
    .ZN(_2262_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _7084_ (.A1(_2261_),
    .A2(_2262_),
    .ZN(_0133_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _7085_ (.A1(_2191_),
    .A2(_2247_),
    .B1(_2250_),
    .B2(\as2650.stack[1][4] ),
    .C(_2244_),
    .ZN(_2263_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _7086_ (.A1(_2186_),
    .A2(_2245_),
    .B(_2263_),
    .ZN(_0134_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _7087_ (.A1(_2197_),
    .A2(_2247_),
    .B1(_2250_),
    .B2(\as2650.stack[1][5] ),
    .C(_2244_),
    .ZN(_2264_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _7088_ (.A1(_2193_),
    .A2(_2245_),
    .B(_2264_),
    .ZN(_0135_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7089_ (.I(_0947_),
    .Z(_2265_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _7090_ (.A1(_2265_),
    .A2(_2247_),
    .B1(_2250_),
    .B2(\as2650.stack[1][6] ),
    .C(_2254_),
    .ZN(_2266_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _7091_ (.A1(_2200_),
    .A2(_2245_),
    .B(_2266_),
    .ZN(_0136_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _7092_ (.A1(_2205_),
    .A2(_2252_),
    .B1(_2253_),
    .B2(\as2650.stack[1][7] ),
    .C(_2243_),
    .ZN(_2267_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _7093_ (.A1(_0951_),
    .A2(_2256_),
    .ZN(_2268_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _7094_ (.A1(_2267_),
    .A2(_2268_),
    .ZN(_0137_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7095_ (.I(\as2650.r123[3][0] ),
    .Z(_2269_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7096_ (.I(_2269_),
    .Z(_0138_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7097_ (.I(\as2650.r123[3][1] ),
    .Z(_2270_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7098_ (.I(_2270_),
    .Z(_0139_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7099_ (.I(\as2650.r123[3][2] ),
    .Z(_2271_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7100_ (.I(_2271_),
    .Z(_0140_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7101_ (.I(\as2650.r123[3][3] ),
    .Z(_2272_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7102_ (.I(_2272_),
    .Z(_0141_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7103_ (.I(\as2650.r123[3][4] ),
    .Z(_2273_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7104_ (.I(_2273_),
    .Z(_0142_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7105_ (.I(\as2650.r123[3][5] ),
    .Z(_2274_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7106_ (.I(_2274_),
    .Z(_0143_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7107_ (.I(\as2650.r123[3][6] ),
    .Z(_2275_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7108_ (.I(_2275_),
    .Z(_0144_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7109_ (.I(\as2650.r123[3][7] ),
    .Z(_2276_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7110_ (.I(_2276_),
    .Z(_0145_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _7111_ (.A1(_0622_),
    .A2(_2208_),
    .ZN(_2277_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7112_ (.I(_2277_),
    .Z(_2278_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7113_ (.I(_2278_),
    .Z(_2279_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _7114_ (.A1(_2148_),
    .A2(_1640_),
    .A3(_2212_),
    .ZN(_2280_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7115_ (.I(_2280_),
    .Z(_2281_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7116_ (.A1(_2165_),
    .A2(_2140_),
    .ZN(_2282_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7117_ (.I(_2282_),
    .Z(_2283_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _7118_ (.A1(_2147_),
    .A2(_2281_),
    .B1(_2283_),
    .B2(\as2650.stack[3][0] ),
    .C(_2278_),
    .ZN(_2284_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _7119_ (.A1(_2138_),
    .A2(_2279_),
    .B(_2284_),
    .ZN(_0146_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7120_ (.I(_0912_),
    .Z(_2285_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7121_ (.I(_2280_),
    .Z(_2286_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7122_ (.I(_2282_),
    .Z(_2287_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7123_ (.I(_2277_),
    .Z(_2288_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _7124_ (.A1(_2285_),
    .A2(_2286_),
    .B1(_2287_),
    .B2(\as2650.stack[3][1] ),
    .C(_2288_),
    .ZN(_2289_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7125_ (.I(_1382_),
    .Z(_2290_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7126_ (.A1(_2215_),
    .A2(_2175_),
    .ZN(_2291_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _7127_ (.A1(_2290_),
    .A2(_2291_),
    .ZN(_2292_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _7128_ (.A1(_2289_),
    .A2(_2292_),
    .ZN(_0147_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _7129_ (.A1(_2258_),
    .A2(_2286_),
    .B1(_2287_),
    .B2(\as2650.stack[3][2] ),
    .C(_2288_),
    .ZN(_2293_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7130_ (.I(_0917_),
    .Z(_2294_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _7131_ (.A1(_2294_),
    .A2(_2291_),
    .ZN(_2295_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _7132_ (.A1(_2293_),
    .A2(_2295_),
    .ZN(_0148_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7133_ (.I(_2182_),
    .Z(_2296_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _7134_ (.A1(_2296_),
    .A2(_2286_),
    .B1(_2287_),
    .B2(\as2650.stack[3][3] ),
    .C(_2288_),
    .ZN(_2297_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7135_ (.I(_0924_),
    .Z(_2298_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _7136_ (.A1(_2298_),
    .A2(_2291_),
    .ZN(_2299_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _7137_ (.A1(_2297_),
    .A2(_2299_),
    .ZN(_0149_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7138_ (.I(_2190_),
    .Z(_2300_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _7139_ (.A1(_2300_),
    .A2(_2281_),
    .B1(_2283_),
    .B2(\as2650.stack[3][4] ),
    .C(_2278_),
    .ZN(_2301_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _7140_ (.A1(_2186_),
    .A2(_2279_),
    .B(_2301_),
    .ZN(_0150_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7141_ (.I(_2196_),
    .Z(_2302_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _7142_ (.A1(_2302_),
    .A2(_2281_),
    .B1(_2283_),
    .B2(\as2650.stack[3][5] ),
    .C(_2278_),
    .ZN(_2303_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _7143_ (.A1(_2193_),
    .A2(_2279_),
    .B(_2303_),
    .ZN(_0151_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _7144_ (.A1(_2265_),
    .A2(_2281_),
    .B1(_2283_),
    .B2(\as2650.stack[3][6] ),
    .C(_2288_),
    .ZN(_2304_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _7145_ (.A1(_2200_),
    .A2(_2279_),
    .B(_2304_),
    .ZN(_0152_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7146_ (.I(_2204_),
    .Z(_2305_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _7147_ (.A1(_2305_),
    .A2(_2286_),
    .B1(_2287_),
    .B2(\as2650.stack[3][7] ),
    .C(_2277_),
    .ZN(_2306_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7148_ (.I(_1411_),
    .Z(_2307_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _7149_ (.A1(_2307_),
    .A2(_2291_),
    .ZN(_2308_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _7150_ (.A1(_2306_),
    .A2(_2308_),
    .ZN(_0153_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _7151_ (.A1(_0857_),
    .A2(_2248_),
    .Z(_2309_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7152_ (.I(_2309_),
    .Z(_2310_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7153_ (.I(_2310_),
    .Z(_2311_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _7154_ (.A1(_0851_),
    .A2(_1921_),
    .A3(_2162_),
    .ZN(_2312_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7155_ (.I(_2312_),
    .Z(_2313_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _7156_ (.A1(_2139_),
    .A2(_1921_),
    .ZN(_2314_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7157_ (.A1(_2165_),
    .A2(_2314_),
    .ZN(_2315_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7158_ (.I(_2315_),
    .Z(_2316_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _7159_ (.A1(_2146_),
    .A2(_2313_),
    .B1(_2316_),
    .B2(\as2650.stack[0][0] ),
    .C(_2310_),
    .ZN(_2317_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _7160_ (.A1(_0848_),
    .A2(_2311_),
    .B(_2317_),
    .ZN(_0154_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7161_ (.I(_2312_),
    .Z(_2318_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7162_ (.I(_2315_),
    .Z(_2319_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7163_ (.I(_2309_),
    .Z(_2320_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _7164_ (.A1(_2285_),
    .A2(_2318_),
    .B1(_2319_),
    .B2(\as2650.stack[0][1] ),
    .C(_2320_),
    .ZN(_2321_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7165_ (.A1(_2175_),
    .A2(_2248_),
    .ZN(_2322_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _7166_ (.A1(_2290_),
    .A2(_2322_),
    .ZN(_2323_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _7167_ (.A1(_2321_),
    .A2(_2323_),
    .ZN(_0155_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _7168_ (.A1(_2258_),
    .A2(_2318_),
    .B1(_2319_),
    .B2(\as2650.stack[0][2] ),
    .C(_2320_),
    .ZN(_2324_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _7169_ (.A1(_2294_),
    .A2(_2322_),
    .ZN(_2325_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _7170_ (.A1(_2324_),
    .A2(_2325_),
    .ZN(_0156_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _7171_ (.A1(_2296_),
    .A2(_2318_),
    .B1(_2319_),
    .B2(\as2650.stack[0][3] ),
    .C(_2320_),
    .ZN(_2326_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _7172_ (.A1(_2298_),
    .A2(_2322_),
    .ZN(_2327_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _7173_ (.A1(_2326_),
    .A2(_2327_),
    .ZN(_0157_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _7174_ (.A1(_2300_),
    .A2(_2313_),
    .B1(_2316_),
    .B2(\as2650.stack[0][4] ),
    .C(_2310_),
    .ZN(_2328_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _7175_ (.A1(_0932_),
    .A2(_2311_),
    .B(_2328_),
    .ZN(_0158_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _7176_ (.A1(_2302_),
    .A2(_2313_),
    .B1(_2316_),
    .B2(\as2650.stack[0][5] ),
    .C(_2310_),
    .ZN(_2329_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _7177_ (.A1(_0938_),
    .A2(_2311_),
    .B(_2329_),
    .ZN(_0159_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _7178_ (.A1(_2265_),
    .A2(_2313_),
    .B1(_2316_),
    .B2(\as2650.stack[0][6] ),
    .C(_2320_),
    .ZN(_2330_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _7179_ (.A1(_2199_),
    .A2(_2311_),
    .B(_2330_),
    .ZN(_0160_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _7180_ (.A1(_2305_),
    .A2(_2318_),
    .B1(_2319_),
    .B2(\as2650.stack[0][7] ),
    .C(_2309_),
    .ZN(_2331_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _7181_ (.A1(_2307_),
    .A2(_2322_),
    .ZN(_2332_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _7182_ (.A1(_2331_),
    .A2(_2332_),
    .ZN(_0161_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _7183_ (.I(\as2650.addr_buff[0] ),
    .ZN(_2333_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _7184_ (.I(_2333_),
    .Z(_2334_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _7185_ (.I(_1272_),
    .Z(_2335_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _7186_ (.I(_1303_),
    .Z(_2336_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7187_ (.A1(_2336_),
    .A2(_4241_),
    .ZN(_2337_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _7188_ (.I(_2337_),
    .Z(_2338_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_2 _7189_ (.A1(_2335_),
    .A2(_2338_),
    .A3(_1324_),
    .A4(_1313_),
    .ZN(_2339_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7190_ (.I(_1338_),
    .Z(_2340_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _7191_ (.A1(_1317_),
    .A2(_2340_),
    .B(_1496_),
    .ZN(_2341_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _7192_ (.A1(_2150_),
    .A2(_1532_),
    .B(_0871_),
    .ZN(_2342_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _7193_ (.A1(_0852_),
    .A2(_1283_),
    .A3(_4253_),
    .ZN(_2343_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_2 _7194_ (.A1(_1351_),
    .A2(_2341_),
    .A3(_2342_),
    .A4(_2343_),
    .ZN(_2344_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _7195_ (.A1(_1086_),
    .A2(_1683_),
    .ZN(_2345_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _7196_ (.A1(_1500_),
    .A2(_1349_),
    .ZN(_2346_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7197_ (.A1(_4393_),
    .A2(_2156_),
    .ZN(_2347_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _7198_ (.I(_0894_),
    .Z(_2348_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _7199_ (.A1(_1464_),
    .A2(_2348_),
    .ZN(_2349_));
 gf180mcu_fd_sc_mcu7t5v0__oai32_1 _7200_ (.A1(_2156_),
    .A2(_1310_),
    .A3(_2346_),
    .B1(_2347_),
    .B2(_2349_),
    .ZN(_2350_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7201_ (.A1(_2345_),
    .A2(_2350_),
    .ZN(_2351_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _7202_ (.A1(_0877_),
    .A2(_1260_),
    .ZN(_2352_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _7203_ (.I(_2352_),
    .Z(_2353_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _7204_ (.I(_1682_),
    .Z(_2354_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _7205_ (.A1(_1524_),
    .A2(_2353_),
    .B(_2354_),
    .ZN(_2355_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _7206_ (.A1(_2351_),
    .A2(_2355_),
    .B(_1701_),
    .ZN(_2356_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_4 _7207_ (.A1(_1569_),
    .A2(_2339_),
    .B(_2344_),
    .C(_2356_),
    .ZN(_2357_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7208_ (.I(_2357_),
    .Z(_2358_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7209_ (.I(_2357_),
    .Z(_2359_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7210_ (.A1(_1691_),
    .A2(_2359_),
    .ZN(_2360_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _7211_ (.A1(_2334_),
    .A2(_2358_),
    .B(_2360_),
    .ZN(_0162_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _7212_ (.I(\as2650.addr_buff[1] ),
    .Z(_2361_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _7213_ (.I(_2361_),
    .Z(_2362_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7214_ (.I(_2357_),
    .Z(_2363_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _7215_ (.A1(_2362_),
    .A2(_2363_),
    .ZN(_2364_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _7216_ (.A1(_1104_),
    .A2(_2358_),
    .B(_2364_),
    .ZN(_0163_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _7217_ (.I(\as2650.addr_buff[2] ),
    .Z(_2365_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _7218_ (.I(_2365_),
    .Z(_2366_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _7219_ (.A1(_2366_),
    .A2(_2363_),
    .ZN(_2367_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _7220_ (.A1(_0376_),
    .A2(_2358_),
    .B(_2367_),
    .ZN(_0164_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _7221_ (.I(\as2650.addr_buff[3] ),
    .ZN(_2368_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7222_ (.I(_2368_),
    .Z(_2369_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7223_ (.I(_2357_),
    .Z(_2370_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7224_ (.A1(_1556_),
    .A2(_2359_),
    .ZN(_2371_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _7225_ (.A1(_2369_),
    .A2(_2370_),
    .B(_2371_),
    .ZN(_0165_));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _7226_ (.I(\as2650.addr_buff[4] ),
    .ZN(_2372_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _7227_ (.I(_1558_),
    .Z(_2373_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7228_ (.A1(_2373_),
    .A2(_2359_),
    .ZN(_2374_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _7229_ (.A1(_2372_),
    .A2(_2370_),
    .B(_2374_),
    .ZN(_0166_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7230_ (.A1(_1292_),
    .A2(_2359_),
    .ZN(_2375_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _7231_ (.A1(_4355_),
    .A2(_2370_),
    .B(_2375_),
    .ZN(_0167_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7232_ (.A1(_1706_),
    .A2(_2363_),
    .ZN(_2376_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _7233_ (.A1(_4357_),
    .A2(_2370_),
    .B(_2376_),
    .ZN(_0168_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _7234_ (.I(_1579_),
    .Z(_2377_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _7235_ (.A1(_1340_),
    .A2(_2363_),
    .ZN(_2378_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _7236_ (.A1(_2377_),
    .A2(_2358_),
    .B(_2378_),
    .ZN(_0169_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _7237_ (.A1(_1309_),
    .A2(_1491_),
    .ZN(_2379_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _7238_ (.A1(_4179_),
    .A2(_1360_),
    .ZN(_2380_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7239_ (.A1(_1252_),
    .A2(_2380_),
    .ZN(_2381_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7240_ (.I(_1479_),
    .Z(_2382_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7241_ (.I(_2382_),
    .Z(_2383_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7242_ (.I(_1489_),
    .Z(_2384_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7243_ (.I(_2384_),
    .Z(_2385_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _7244_ (.I(_2385_),
    .Z(_2386_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7245_ (.I(_1466_),
    .Z(_2387_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7246_ (.I(_2387_),
    .Z(_2388_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _7247_ (.A1(_2383_),
    .A2(_2386_),
    .A3(_2380_),
    .A4(_2388_),
    .ZN(_2389_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _7248_ (.A1(_1367_),
    .A2(_1279_),
    .A3(_2346_),
    .ZN(_2390_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7249_ (.I(_1321_),
    .Z(_2391_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _7250_ (.A1(_1486_),
    .A2(_2391_),
    .A3(_1702_),
    .ZN(_2392_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _7251_ (.A1(_2381_),
    .A2(_2389_),
    .A3(_2390_),
    .A4(_2392_),
    .ZN(_2393_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _7252_ (.A1(_1366_),
    .A2(_2379_),
    .A3(_2393_),
    .ZN(_2394_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _7253_ (.I(_4176_),
    .Z(_2395_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _7254_ (.I(_2395_),
    .Z(_2396_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _7255_ (.A1(_1451_),
    .A2(_2396_),
    .B(_1350_),
    .ZN(_2397_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _7256_ (.A1(net24),
    .A2(_2394_),
    .ZN(_2398_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _7257_ (.A1(_2394_),
    .A2(_2397_),
    .B(_2398_),
    .C(_1410_),
    .ZN(_0170_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _7258_ (.I(_1571_),
    .Z(_2399_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _7259_ (.A1(_1319_),
    .A2(_1347_),
    .ZN(_2400_));
 gf180mcu_fd_sc_mcu7t5v0__and4_1 _7260_ (.A1(_2399_),
    .A2(_1278_),
    .A3(_1242_),
    .A4(_2400_),
    .Z(_2401_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _7261_ (.A1(net22),
    .A2(_2401_),
    .ZN(_2402_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _7262_ (.A1(_4323_),
    .A2(_2401_),
    .B(_2402_),
    .C(_1410_),
    .ZN(_0171_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _7263_ (.I(_1327_),
    .Z(_2403_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7264_ (.A1(_1282_),
    .A2(_1361_),
    .ZN(_2404_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _7265_ (.A1(_2383_),
    .A2(_1547_),
    .B(_2404_),
    .ZN(_2405_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _7266_ (.I(_1325_),
    .Z(_2406_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _7267_ (.I(_2406_),
    .Z(_2407_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _7268_ (.I(_1321_),
    .Z(_2408_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _7269_ (.A1(_1260_),
    .A2(_1248_),
    .ZN(_2409_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _7270_ (.I(_0896_),
    .Z(_2410_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_4 _7271_ (.A1(_1356_),
    .A2(_1513_),
    .A3(_2410_),
    .A4(_1370_),
    .ZN(_2411_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_4 _7272_ (.A1(_2407_),
    .A2(_2408_),
    .B1(_1483_),
    .B2(_2409_),
    .C(_2411_),
    .ZN(_2412_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_2 _7273_ (.A1(_2403_),
    .A2(_2405_),
    .B(_2412_),
    .C(_2400_),
    .ZN(_2413_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7274_ (.A1(net23),
    .A2(_2413_),
    .ZN(_2414_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _7275_ (.A1(_4209_),
    .A2(_2413_),
    .B(_2414_),
    .C(_1566_),
    .ZN(_0172_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7276_ (.I(_1301_),
    .Z(_2415_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _7277_ (.I(_2415_),
    .Z(_2416_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7278_ (.I(net28),
    .Z(_2417_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7279_ (.I(_2417_),
    .Z(_2418_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _7280_ (.A1(_4199_),
    .A2(_4544_),
    .ZN(_2419_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_2 _7281_ (.A1(_0654_),
    .A2(_1493_),
    .A3(_2419_),
    .ZN(_2420_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _7282_ (.A1(_4551_),
    .A2(_1501_),
    .ZN(_2421_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7283_ (.A1(_2420_),
    .A2(_2421_),
    .ZN(_2422_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _7284_ (.A1(_4427_),
    .A2(_1240_),
    .A3(_4425_),
    .ZN(_2423_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_1 _7285_ (.A1(_0654_),
    .A2(_1253_),
    .A3(_1468_),
    .B(_2423_),
    .ZN(_2424_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _7286_ (.A1(_2419_),
    .A2(_2424_),
    .B(_4418_),
    .ZN(_2425_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7287_ (.A1(_2422_),
    .A2(_2425_),
    .ZN(_2426_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _7288_ (.A1(_1471_),
    .A2(_1501_),
    .ZN(_2427_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _7289_ (.A1(_1230_),
    .A2(_2427_),
    .B(_1350_),
    .ZN(_2428_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _7290_ (.A1(_1095_),
    .A2(_1324_),
    .ZN(_2429_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _7291_ (.A1(_1939_),
    .A2(_2429_),
    .A3(_1347_),
    .ZN(_2430_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _7292_ (.A1(_1163_),
    .A2(_2408_),
    .B(_2406_),
    .ZN(_2431_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7293_ (.A1(_4169_),
    .A2(_4237_),
    .ZN(_2432_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7294_ (.A1(_1355_),
    .A2(_2432_),
    .ZN(_2433_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7295_ (.A1(_1312_),
    .A2(_2433_),
    .ZN(_2434_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _7296_ (.A1(_4233_),
    .A2(_1326_),
    .A3(_2434_),
    .ZN(_2435_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7297_ (.A1(_1314_),
    .A2(_2435_),
    .ZN(_2436_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _7298_ (.A1(_1497_),
    .A2(_4543_),
    .ZN(_2437_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _7299_ (.I(_0869_),
    .Z(_2438_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _7300_ (.A1(_4423_),
    .A2(_1257_),
    .Z(_2439_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _7301_ (.A1(_4431_),
    .A2(_1256_),
    .B(_2439_),
    .ZN(_2440_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _7302_ (.A1(_2437_),
    .A2(_2438_),
    .A3(_2440_),
    .ZN(_2441_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _7303_ (.A1(_4200_),
    .A2(_1364_),
    .A3(_1363_),
    .ZN(_2442_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _7304_ (.A1(_1497_),
    .A2(_4250_),
    .ZN(_2443_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _7305_ (.A1(_1346_),
    .A2(_1683_),
    .A3(_2443_),
    .ZN(_2444_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_2 _7306_ (.A1(_2436_),
    .A2(_2441_),
    .A3(_2442_),
    .A4(_2444_),
    .ZN(_2445_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_2 _7307_ (.A1(_4422_),
    .A2(_4430_),
    .A3(_4432_),
    .A4(_1470_),
    .ZN(_2446_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7308_ (.A1(_1087_),
    .A2(_2446_),
    .ZN(_2447_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_4 _7309_ (.A1(_1230_),
    .A2(_1471_),
    .A3(_1231_),
    .A4(_1368_),
    .ZN(_2448_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _7310_ (.A1(_0469_),
    .A2(_1261_),
    .A3(_4425_),
    .ZN(_2449_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _7311_ (.A1(_4442_),
    .A2(_2449_),
    .Z(_2450_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _7312_ (.A1(_4220_),
    .A2(_2406_),
    .B(_0970_),
    .ZN(_2451_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _7313_ (.A1(_2450_),
    .A2(_1503_),
    .A3(_2451_),
    .ZN(_2452_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _7314_ (.A1(_2406_),
    .A2(_2448_),
    .B(_2452_),
    .ZN(_2453_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_1 _7315_ (.A1(_1501_),
    .A2(_1504_),
    .A3(_2351_),
    .B(_2453_),
    .ZN(_2454_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _7316_ (.A1(_2445_),
    .A2(_2447_),
    .A3(_2454_),
    .ZN(_2455_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _7317_ (.A1(_2428_),
    .A2(_2430_),
    .A3(_2431_),
    .A4(_2455_),
    .ZN(_2456_));
 gf180mcu_fd_sc_mcu7t5v0__or4_1 _7318_ (.A1(_1316_),
    .A2(_4443_),
    .A3(_0397_),
    .A4(_0339_),
    .Z(_2457_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_2 _7319_ (.A1(_0717_),
    .A2(_0762_),
    .Z(_2458_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_2 _7320_ (.A1(_4398_),
    .A2(_1106_),
    .A3(_0378_),
    .ZN(_2459_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_4 _7321_ (.A1(_0512_),
    .A2(_0603_),
    .A3(_0690_),
    .A4(_2459_),
    .ZN(_2460_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_4 _7322_ (.A1(_4161_),
    .A2(_2458_),
    .A3(_0833_),
    .A4(_2460_),
    .ZN(_2461_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _7323_ (.A1(_2437_),
    .A2(_2438_),
    .A3(_2461_),
    .ZN(_2462_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7324_ (.A1(_2457_),
    .A2(_2462_),
    .ZN(_2463_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _7325_ (.A1(_2426_),
    .A2(_2456_),
    .A3(_2463_),
    .ZN(_2464_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7326_ (.I(_2464_),
    .Z(_2465_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7327_ (.I(_2465_),
    .Z(_2466_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7328_ (.I(_1308_),
    .Z(_2467_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7329_ (.A1(_4349_),
    .A2(_4347_),
    .ZN(_2468_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7330_ (.I(_2468_),
    .Z(_2469_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7331_ (.A1(_2469_),
    .A2(_4352_),
    .ZN(_2470_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _7332_ (.A1(_1550_),
    .A2(_2470_),
    .Z(_2471_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7333_ (.I(_4267_),
    .Z(_2472_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7334_ (.I(_2472_),
    .Z(_2473_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7335_ (.A1(_2473_),
    .A2(_4361_),
    .ZN(_2474_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _7336_ (.A1(_1550_),
    .A2(_2474_),
    .Z(_2475_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7337_ (.I(_1341_),
    .Z(_2476_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7338_ (.I(_2476_),
    .Z(_2477_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _7339_ (.A1(_2467_),
    .A2(_2471_),
    .B1(_2475_),
    .B2(_2477_),
    .ZN(_2478_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_2 _7340_ (.A1(_1678_),
    .A2(_1676_),
    .A3(_4240_),
    .ZN(_2479_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7341_ (.I(_2479_),
    .Z(_2480_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7342_ (.I(_0853_),
    .Z(_2481_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _7343_ (.I(_2481_),
    .Z(_2482_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7344_ (.A1(_1463_),
    .A2(_2482_),
    .ZN(_2483_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _7345_ (.I(_0885_),
    .Z(_2484_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7346_ (.A1(_2484_),
    .A2(_1311_),
    .ZN(_2485_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7347_ (.I(_2485_),
    .Z(_2486_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _7348_ (.A1(_0863_),
    .A2(_4391_),
    .Z(_2487_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _7349_ (.A1(_2486_),
    .A2(_2487_),
    .ZN(_2488_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _7350_ (.A1(_2418_),
    .A2(_2480_),
    .B(_2483_),
    .C(_2488_),
    .ZN(_2489_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _7351_ (.A1(_1311_),
    .A2(_2478_),
    .B(_2489_),
    .ZN(_2490_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7352_ (.A1(_1482_),
    .A2(_2481_),
    .ZN(_2491_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7353_ (.I(_2491_),
    .Z(_2492_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _7354_ (.A1(_2150_),
    .A2(_4393_),
    .ZN(_2493_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7355_ (.I(_2493_),
    .Z(_2494_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7356_ (.I(_2494_),
    .Z(_2495_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _7357_ (.A1(_2492_),
    .A2(_2495_),
    .ZN(_2496_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7358_ (.A1(_1545_),
    .A2(_2487_),
    .ZN(_2497_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _7359_ (.A1(_2418_),
    .A2(_1710_),
    .B(_2497_),
    .ZN(_2498_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7360_ (.A1(_0872_),
    .A2(_2151_),
    .ZN(_2499_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7361_ (.I(_2499_),
    .Z(_2500_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _7362_ (.A1(_2396_),
    .A2(_1684_),
    .ZN(_2501_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7363_ (.I(_2501_),
    .Z(_2502_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _7364_ (.I(_0882_),
    .Z(_2503_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _7365_ (.A1(_2153_),
    .A2(_2503_),
    .ZN(_2504_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7366_ (.I(_2504_),
    .Z(_2505_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _7367_ (.A1(_0881_),
    .A2(_2154_),
    .Z(_2506_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7368_ (.I(_2506_),
    .Z(_2507_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7369_ (.I(_2507_),
    .Z(_2508_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _7370_ (.I(_2410_),
    .Z(_2509_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _7371_ (.A1(_2417_),
    .A2(_2509_),
    .ZN(_2510_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _7372_ (.A1(_2418_),
    .A2(_2505_),
    .B1(_2508_),
    .B2(_1551_),
    .C(_2510_),
    .ZN(_2511_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _7373_ (.A1(_2498_),
    .A2(_2500_),
    .B1(_2502_),
    .B2(_2511_),
    .ZN(_2512_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7374_ (.I(_2492_),
    .Z(_2513_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _7375_ (.I(_1374_),
    .Z(_2514_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_1 _7376_ (.A1(_2145_),
    .A2(_2496_),
    .B1(_2512_),
    .B2(_2513_),
    .C(_2514_),
    .ZN(_2515_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _7377_ (.A1(_2490_),
    .A2(_2515_),
    .B(_2403_),
    .ZN(_2516_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7378_ (.I(_1359_),
    .Z(_2517_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _7379_ (.A1(_0865_),
    .A2(_2517_),
    .B(_2465_),
    .ZN(_2518_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _7380_ (.A1(_2418_),
    .A2(_2466_),
    .B1(_2516_),
    .B2(_2518_),
    .ZN(_2519_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _7381_ (.A1(_2416_),
    .A2(_2519_),
    .ZN(_0173_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7382_ (.I(_2464_),
    .Z(_2520_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7383_ (.I(_2520_),
    .Z(_2521_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7384_ (.I(_2517_),
    .Z(_2522_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _7385_ (.A1(_1498_),
    .A2(_4418_),
    .ZN(_2523_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7386_ (.I(_2523_),
    .Z(_2524_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _7387_ (.I(_2524_),
    .Z(_2525_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7388_ (.A1(_1695_),
    .A2(_2395_),
    .ZN(_2526_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7389_ (.I(_2526_),
    .Z(_2527_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7390_ (.A1(_2525_),
    .A2(_2527_),
    .ZN(_2528_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7391_ (.A1(_1260_),
    .A2(_0872_),
    .ZN(_2529_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _7392_ (.I(net29),
    .Z(_2530_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _7393_ (.A1(_2153_),
    .A2(_2384_),
    .Z(_2531_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7394_ (.I(_2531_),
    .Z(_2532_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _7395_ (.I(_0896_),
    .Z(_2533_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7396_ (.A1(_1340_),
    .A2(_2533_),
    .ZN(_2534_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _7397_ (.I(_2534_),
    .Z(_2535_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _7398_ (.I(_4531_),
    .Z(_2536_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _7399_ (.A1(_2530_),
    .A2(_2417_),
    .Z(_2537_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _7400_ (.I(_2154_),
    .Z(_2538_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _7401_ (.I(_2538_),
    .Z(_2539_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7402_ (.I(_2539_),
    .Z(_2540_));
 gf180mcu_fd_sc_mcu7t5v0__oai222_1 _7403_ (.A1(_2530_),
    .A2(_2532_),
    .B1(_2535_),
    .B2(_2536_),
    .C1(_2537_),
    .C2(_2540_),
    .ZN(_2541_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7404_ (.I(_1336_),
    .Z(_2542_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7405_ (.A1(\as2650.pc[0] ),
    .A2(net6),
    .ZN(_2543_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _7406_ (.A1(_0910_),
    .A2(_4528_),
    .Z(_2544_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _7407_ (.A1(_2543_),
    .A2(_2544_),
    .Z(_2545_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7408_ (.A1(_2542_),
    .A2(_2545_),
    .ZN(_2546_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _7409_ (.A1(_2530_),
    .A2(_1619_),
    .B(_2499_),
    .C(_2546_),
    .ZN(_2547_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _7410_ (.A1(_2529_),
    .A2(_2541_),
    .B(_2547_),
    .ZN(_2548_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7411_ (.I(_2523_),
    .Z(_2549_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7412_ (.I(_2549_),
    .Z(_2550_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _7413_ (.I(_1569_),
    .Z(_2551_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _7414_ (.A1(_0911_),
    .A2(_2528_),
    .B1(_2548_),
    .B2(_2550_),
    .C(_2551_),
    .ZN(_2552_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7415_ (.I(_2469_),
    .Z(_2553_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7416_ (.I(_1308_),
    .Z(_2554_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7417_ (.I(_2468_),
    .Z(_2555_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7418_ (.A1(_4390_),
    .A2(_4352_),
    .ZN(_2556_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _7419_ (.A1(_4529_),
    .A2(_0292_),
    .A3(_2556_),
    .Z(_2557_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7420_ (.A1(_2555_),
    .A2(_2557_),
    .ZN(_2558_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _7421_ (.A1(_2536_),
    .A2(_2553_),
    .B(_2554_),
    .C(_2558_),
    .ZN(_2559_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7422_ (.I(_2472_),
    .Z(_2560_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7423_ (.A1(_4390_),
    .A2(_4360_),
    .ZN(_2561_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _7424_ (.A1(_4529_),
    .A2(_4513_),
    .A3(_2561_),
    .Z(_2562_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7425_ (.A1(_2473_),
    .A2(_2562_),
    .ZN(_2563_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7426_ (.I(_1341_),
    .Z(_2564_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7427_ (.I(_2564_),
    .Z(_2565_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _7428_ (.A1(_2536_),
    .A2(_2560_),
    .B(_2563_),
    .C(_2565_),
    .ZN(_2566_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7429_ (.A1(_2559_),
    .A2(_2566_),
    .ZN(_2567_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _7430_ (.A1(_0862_),
    .A2(_4390_),
    .ZN(_2568_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _7431_ (.A1(_2568_),
    .A2(_2544_),
    .Z(_2569_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7432_ (.I(_1344_),
    .Z(_2570_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _7433_ (.A1(_2486_),
    .A2(_2569_),
    .B(_2570_),
    .ZN(_2571_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _7434_ (.A1(_2480_),
    .A2(_2537_),
    .B1(_2567_),
    .B2(_1337_),
    .C(_2571_),
    .ZN(_2572_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7435_ (.I(_1357_),
    .Z(_2573_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _7436_ (.A1(_2552_),
    .A2(_2572_),
    .B(_2573_),
    .ZN(_2574_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _7437_ (.A1(_0912_),
    .A2(_2522_),
    .B(_2574_),
    .ZN(_2575_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _7438_ (.A1(_2530_),
    .A2(_2520_),
    .ZN(_2576_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7439_ (.I(_1390_),
    .Z(_2577_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _7440_ (.I(_2577_),
    .Z(_2578_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _7441_ (.A1(_2521_),
    .A2(_2575_),
    .B(_2576_),
    .C(_2578_),
    .ZN(_0174_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7442_ (.I(_2520_),
    .Z(_2579_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7443_ (.I(_2517_),
    .Z(_2580_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7444_ (.I(net7),
    .Z(_2581_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _7445_ (.A1(_0289_),
    .A2(_0291_),
    .B(_2581_),
    .ZN(_2582_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _7446_ (.A1(_2581_),
    .A2(_0289_),
    .A3(_0291_),
    .ZN(_2583_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _7447_ (.A1(_2556_),
    .A2(_2582_),
    .B(_2583_),
    .ZN(_2584_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _7448_ (.A1(_0351_),
    .A2(_0357_),
    .B(_0374_),
    .ZN(_2585_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7449_ (.A1(_1554_),
    .A2(_0358_),
    .ZN(_2586_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7450_ (.A1(_2585_),
    .A2(_2586_),
    .ZN(_2587_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7451_ (.I(_4246_),
    .Z(_2588_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _7452_ (.A1(_2584_),
    .A2(_2587_),
    .B(_2588_),
    .ZN(_2589_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _7453_ (.A1(_2584_),
    .A2(_2587_),
    .B(_2589_),
    .ZN(_2590_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _7454_ (.A1(_1699_),
    .A2(_2553_),
    .B(_2467_),
    .C(_2590_),
    .ZN(_2591_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_4 _7455_ (.A1(_4503_),
    .A2(_0350_),
    .B1(_0356_),
    .B2(_0386_),
    .C(_0387_),
    .ZN(_2592_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _7456_ (.A1(_4511_),
    .A2(_4512_),
    .B(_4528_),
    .ZN(_2593_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _7457_ (.A1(_4528_),
    .A2(_4511_),
    .A3(_4512_),
    .ZN(_2594_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _7458_ (.A1(_2593_),
    .A2(_2561_),
    .B(_2594_),
    .ZN(_2595_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _7459_ (.A1(_1553_),
    .A2(_2592_),
    .A3(_2595_),
    .Z(_2596_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7460_ (.A1(_2560_),
    .A2(_2596_),
    .ZN(_2597_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7461_ (.I(_2564_),
    .Z(_2598_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _7462_ (.A1(_1555_),
    .A2(_2560_),
    .B(_2597_),
    .C(_2598_),
    .ZN(_2599_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7463_ (.A1(_2591_),
    .A2(_2599_),
    .ZN(_2600_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _7464_ (.A1(\as2650.pc[2] ),
    .A2(net8),
    .Z(_2601_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7465_ (.I(_2601_),
    .Z(_2602_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _7466_ (.A1(\as2650.pc[1] ),
    .A2(net7),
    .ZN(_2603_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7467_ (.A1(_0909_),
    .A2(net7),
    .ZN(_2604_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _7468_ (.A1(_2568_),
    .A2(_2603_),
    .B(_2604_),
    .ZN(_2605_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _7469_ (.A1(_2602_),
    .A2(_2605_),
    .Z(_2606_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _7470_ (.I(_1338_),
    .Z(_2607_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _7471_ (.A1(_2602_),
    .A2(_2605_),
    .B(_2607_),
    .ZN(_2608_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _7472_ (.I(net30),
    .Z(_2609_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7473_ (.A1(net29),
    .A2(_2417_),
    .ZN(_2610_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _7474_ (.A1(_2609_),
    .A2(_2610_),
    .Z(_2611_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7475_ (.I(_1306_),
    .Z(_2612_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _7476_ (.I(_2612_),
    .Z(_2613_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_1 _7477_ (.A1(_2606_),
    .A2(_2608_),
    .B1(_2611_),
    .B2(_2613_),
    .C(_2570_),
    .ZN(_2614_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _7478_ (.A1(_1337_),
    .A2(_2600_),
    .B(_2614_),
    .ZN(_2615_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _7479_ (.A1(_2540_),
    .A2(_2611_),
    .ZN(_2616_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _7480_ (.A1(_2609_),
    .A2(_2505_),
    .B1(_2508_),
    .B2(_1555_),
    .C(_2616_),
    .ZN(_2617_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _7481_ (.I(_2542_),
    .Z(_2618_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _7482_ (.A1(_2543_),
    .A2(_2603_),
    .B(_2604_),
    .ZN(_2619_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _7483_ (.A1(_2602_),
    .A2(_2619_),
    .ZN(_2620_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7484_ (.A1(_1545_),
    .A2(_2620_),
    .ZN(_2621_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _7485_ (.A1(_2609_),
    .A2(_2618_),
    .B(_2500_),
    .C(_2621_),
    .ZN(_2622_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _7486_ (.A1(_2529_),
    .A2(_2617_),
    .B(_2622_),
    .ZN(_2623_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _7487_ (.I(_1569_),
    .Z(_2624_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _7488_ (.A1(_0921_),
    .A2(_2528_),
    .B1(_2623_),
    .B2(_2550_),
    .C(_2624_),
    .ZN(_2625_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _7489_ (.A1(_2615_),
    .A2(_2625_),
    .B(_2573_),
    .ZN(_2626_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _7490_ (.A1(_2178_),
    .A2(_2580_),
    .B(_2626_),
    .ZN(_2627_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _7491_ (.A1(_2609_),
    .A2(_2466_),
    .B(_1635_),
    .ZN(_2628_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _7492_ (.A1(_2579_),
    .A2(_2627_),
    .B(_2628_),
    .ZN(_0175_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7493_ (.I(_1283_),
    .Z(_2629_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _7494_ (.I(_2629_),
    .Z(_2630_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7495_ (.I(_2443_),
    .Z(_2631_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _7496_ (.I(_2631_),
    .Z(_2632_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _7497_ (.I(_2632_),
    .Z(_2633_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7498_ (.I(_1532_),
    .Z(_2634_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _7499_ (.I(_2634_),
    .Z(_2635_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _7500_ (.A1(_2181_),
    .A2(_0506_),
    .ZN(_2636_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _7501_ (.A1(_0926_),
    .A2(_1584_),
    .ZN(_2637_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _7502_ (.A1(_2636_),
    .A2(_2637_),
    .ZN(_2638_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _7503_ (.A1(\as2650.pc[2] ),
    .A2(_0373_),
    .Z(_2639_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _7504_ (.A1(_2602_),
    .A2(_2619_),
    .B(_2639_),
    .ZN(_2640_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _7505_ (.A1(_2638_),
    .A2(_2640_),
    .Z(_2641_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _7506_ (.A1(_1614_),
    .A2(_2641_),
    .Z(_2642_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _7507_ (.I(net31),
    .Z(_2643_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7508_ (.I(_1579_),
    .Z(_2644_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7509_ (.I(_2352_),
    .Z(_2645_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _7510_ (.A1(_1684_),
    .A2(_2645_),
    .ZN(_2646_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _7511_ (.A1(_2643_),
    .A2(_2644_),
    .B(_2646_),
    .ZN(_2647_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _7512_ (.I(_2384_),
    .Z(_2648_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _7513_ (.A1(net30),
    .A2(net29),
    .A3(net28),
    .ZN(_2649_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _7514_ (.A1(_2643_),
    .A2(_2649_),
    .Z(_2650_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _7515_ (.A1(_0508_),
    .A2(_1489_),
    .ZN(_2651_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _7516_ (.A1(_2648_),
    .A2(_2650_),
    .B1(_2651_),
    .B2(_1340_),
    .ZN(_2652_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _7517_ (.A1(_2643_),
    .A2(_2532_),
    .B(_2652_),
    .ZN(_2653_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _7518_ (.A1(_2642_),
    .A2(_2647_),
    .B1(_2653_),
    .B2(_2502_),
    .ZN(_2654_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7519_ (.A1(_2335_),
    .A2(_2527_),
    .ZN(_2655_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7520_ (.A1(_0928_),
    .A2(_2655_),
    .ZN(_2656_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _7521_ (.A1(_2635_),
    .A2(_2654_),
    .B(_2656_),
    .ZN(_2657_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _7522_ (.I(_2340_),
    .Z(_2658_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _7523_ (.A1(_2639_),
    .A2(_2606_),
    .ZN(_2659_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _7524_ (.A1(_2638_),
    .A2(_2659_),
    .ZN(_2660_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7525_ (.A1(_2336_),
    .A2(_2479_),
    .ZN(_2661_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7526_ (.I(_1308_),
    .Z(_2662_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _7527_ (.A1(_1585_),
    .A2(_0485_),
    .Z(_2663_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _7528_ (.A1(_1584_),
    .A2(_0479_),
    .A3(_0484_),
    .ZN(_2664_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _7529_ (.A1(_2663_),
    .A2(_2664_),
    .ZN(_2665_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_2 _7530_ (.A1(_0374_),
    .A2(_0351_),
    .A3(_0357_),
    .ZN(_2666_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _7531_ (.A1(_2584_),
    .A2(_2585_),
    .B(_2666_),
    .ZN(_2667_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _7532_ (.A1(_2665_),
    .A2(_2667_),
    .ZN(_2668_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7533_ (.A1(_2469_),
    .A2(_2668_),
    .ZN(_2669_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _7534_ (.A1(_1594_),
    .A2(_2555_),
    .B(_2662_),
    .C(_2669_),
    .ZN(_2670_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7535_ (.A1(_0375_),
    .A2(_2592_),
    .ZN(_2671_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_2 _7536_ (.A1(_0374_),
    .A2(_2592_),
    .B1(_2593_),
    .B2(_2561_),
    .C(_2594_),
    .ZN(_2672_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7537_ (.A1(_2671_),
    .A2(_2672_),
    .ZN(_2673_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _7538_ (.A1(_1585_),
    .A2(_0491_),
    .A3(_2673_),
    .Z(_2674_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7539_ (.A1(_2472_),
    .A2(_2674_),
    .ZN(_2675_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _7540_ (.A1(_1594_),
    .A2(_2473_),
    .B(_2675_),
    .C(_2564_),
    .ZN(_2676_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7541_ (.A1(_2670_),
    .A2(_2676_),
    .ZN(_2677_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _7542_ (.A1(_2661_),
    .A2(_2677_),
    .B1(_2650_),
    .B2(_2479_),
    .C(_2340_),
    .ZN(_2678_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _7543_ (.A1(_2658_),
    .A2(_2660_),
    .B(_2678_),
    .C(_2483_),
    .ZN(_2679_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _7544_ (.A1(_0928_),
    .A2(_2630_),
    .B1(_2633_),
    .B2(_2657_),
    .C(_2679_),
    .ZN(_2680_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7545_ (.I(_2403_),
    .Z(_2681_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _7546_ (.A1(_2183_),
    .A2(_2580_),
    .B1(_2680_),
    .B2(_2681_),
    .ZN(_2682_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _7547_ (.A1(_2643_),
    .A2(_2466_),
    .B(_1635_),
    .ZN(_2683_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _7548_ (.A1(_2579_),
    .A2(_2682_),
    .B(_2683_),
    .ZN(_0176_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7549_ (.I(_2517_),
    .Z(_2684_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7550_ (.A1(_2190_),
    .A2(_2655_),
    .ZN(_2685_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _7551_ (.I(_1513_),
    .Z(_2686_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _7552_ (.I(net32),
    .Z(_2687_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7553_ (.I(_2507_),
    .Z(_2688_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _7554_ (.I(net31),
    .ZN(_2689_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _7555_ (.A1(_2689_),
    .A2(_2649_),
    .ZN(_2690_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _7556_ (.A1(_2687_),
    .A2(_2690_),
    .ZN(_2691_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _7557_ (.A1(_1582_),
    .A2(_2688_),
    .B1(_2691_),
    .B2(_2648_),
    .ZN(_2692_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _7558_ (.A1(_2687_),
    .A2(_2532_),
    .B(_2502_),
    .C(_2692_),
    .ZN(_2693_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7559_ (.I(_0594_),
    .Z(_2694_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _7560_ (.A1(_2187_),
    .A2(_2694_),
    .Z(_2695_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _7561_ (.A1(_2601_),
    .A2(_2619_),
    .B(_2637_),
    .C(_2639_),
    .ZN(_2696_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _7562_ (.A1(_2636_),
    .A2(_2696_),
    .Z(_2697_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _7563_ (.A1(_2695_),
    .A2(_2697_),
    .Z(_2698_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7564_ (.A1(_1545_),
    .A2(_2698_),
    .ZN(_2699_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _7565_ (.A1(_2687_),
    .A2(_1710_),
    .B(_2500_),
    .C(_2699_),
    .ZN(_2700_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _7566_ (.A1(_2693_),
    .A2(_2700_),
    .B(_1252_),
    .ZN(_2701_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _7567_ (.A1(_2190_),
    .A2(_2686_),
    .B1(_1701_),
    .B2(_2701_),
    .ZN(_2702_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _7568_ (.A1(\as2650.addr_buff[7] ),
    .A2(_4266_),
    .Z(_2703_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7569_ (.I(_2703_),
    .Z(_2704_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7570_ (.A1(_2565_),
    .A2(_2704_),
    .ZN(_2705_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _7571_ (.A1(_0507_),
    .A2(_0490_),
    .ZN(_2706_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_2 _7572_ (.A1(_0507_),
    .A2(_0490_),
    .B1(_2671_),
    .B2(_2672_),
    .ZN(_2707_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _7573_ (.A1(_2706_),
    .A2(_2707_),
    .ZN(_2708_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _7574_ (.A1(_1581_),
    .A2(_0578_),
    .A3(_2708_),
    .Z(_2709_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_2 _7575_ (.A1(_2584_),
    .A2(_2585_),
    .B(_2666_),
    .C(_2664_),
    .ZN(_2710_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _7576_ (.A1(_2663_),
    .A2(_2710_),
    .ZN(_2711_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _7577_ (.A1(_1580_),
    .A2(_0614_),
    .A3(_2711_),
    .Z(_2712_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7578_ (.A1(_2555_),
    .A2(_2712_),
    .ZN(_2713_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _7579_ (.A1(_0597_),
    .A2(_2553_),
    .B(_2554_),
    .C(_2713_),
    .ZN(_2714_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_1 _7580_ (.A1(_1582_),
    .A2(_2705_),
    .B1(_2709_),
    .B2(_4268_),
    .C(_2714_),
    .ZN(_2715_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7581_ (.A1(_2181_),
    .A2(_0507_),
    .ZN(_2716_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _7582_ (.A1(_2636_),
    .A2(_2659_),
    .B(_2716_),
    .ZN(_2717_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _7583_ (.A1(_2695_),
    .A2(_2717_),
    .Z(_2718_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _7584_ (.I(_2340_),
    .Z(_2719_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _7585_ (.I(_2612_),
    .Z(_2720_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _7586_ (.A1(_2720_),
    .A2(_2691_),
    .B(_2570_),
    .ZN(_2721_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _7587_ (.A1(_1337_),
    .A2(_2715_),
    .B1(_2718_),
    .B2(_2719_),
    .C(_2721_),
    .ZN(_2722_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _7588_ (.A1(_2685_),
    .A2(_2702_),
    .B(_2722_),
    .ZN(_2723_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _7589_ (.A1(_2191_),
    .A2(_2684_),
    .B1(_2723_),
    .B2(_2681_),
    .ZN(_2724_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _7590_ (.A1(_2687_),
    .A2(_2466_),
    .B(_1635_),
    .ZN(_2725_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _7591_ (.A1(_2579_),
    .A2(_2724_),
    .B(_2725_),
    .ZN(_0177_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _7592_ (.A1(_0939_),
    .A2(net1),
    .Z(_2726_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _7593_ (.I(_2726_),
    .Z(_2727_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7594_ (.A1(_2188_),
    .A2(_0596_),
    .ZN(_2728_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7595_ (.A1(_2695_),
    .A2(_2717_),
    .ZN(_2729_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7596_ (.A1(_2728_),
    .A2(_2729_),
    .ZN(_2730_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _7597_ (.A1(_2727_),
    .A2(_2730_),
    .ZN(_2731_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _7598_ (.A1(_0594_),
    .A2(_0613_),
    .ZN(_2732_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7599_ (.A1(_2694_),
    .A2(_0613_),
    .ZN(_2733_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_2 _7600_ (.A1(_2663_),
    .A2(_2732_),
    .A3(_2710_),
    .B(_2733_),
    .ZN(_2734_));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_1 _7601_ (.A1(_1180_),
    .A2(_0668_),
    .A3(_2734_),
    .ZN(_2735_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _7602_ (.I(_0684_),
    .Z(_2736_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7603_ (.A1(_2736_),
    .A2(_4246_),
    .ZN(_2737_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _7604_ (.A1(_2588_),
    .A2(_2735_),
    .B(_2737_),
    .C(_2662_),
    .ZN(_2738_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _7605_ (.A1(_0595_),
    .A2(_0577_),
    .ZN(_2739_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7606_ (.A1(_0595_),
    .A2(_0577_),
    .ZN(_2740_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_2 _7607_ (.A1(_2706_),
    .A2(_2739_),
    .A3(_2707_),
    .B(_2740_),
    .ZN(_2741_));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_1 _7608_ (.A1(_1180_),
    .A2(_0698_),
    .A3(_2741_),
    .ZN(_2742_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7609_ (.A1(_0685_),
    .A2(_2703_),
    .ZN(_2743_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7610_ (.I(_1341_),
    .Z(_2744_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _7611_ (.A1(_2704_),
    .A2(_2742_),
    .B(_2743_),
    .C(_2744_),
    .ZN(_2745_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7612_ (.A1(_2738_),
    .A2(_2745_),
    .ZN(_2746_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _7613_ (.A1(net32),
    .A2(_2690_),
    .Z(_2747_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _7614_ (.A1(net33),
    .A2(_2747_),
    .Z(_2748_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _7615_ (.I(_2748_),
    .ZN(_2749_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _7616_ (.A1(_2661_),
    .A2(_2746_),
    .B1(_2749_),
    .B2(_2480_),
    .C(_2658_),
    .ZN(_2750_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7617_ (.I(_2483_),
    .Z(_2751_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _7618_ (.A1(_2719_),
    .A2(_2731_),
    .B(_2750_),
    .C(_2751_),
    .ZN(_2752_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _7619_ (.I(_1701_),
    .Z(_2753_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7620_ (.I(_2154_),
    .Z(_2754_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _7621_ (.I(_2754_),
    .Z(_2755_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _7622_ (.I(_2755_),
    .Z(_2756_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7623_ (.I(net33),
    .Z(_2757_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _7624_ (.A1(_2757_),
    .A2(_2504_),
    .B1(_2688_),
    .B2(_2736_),
    .C(_2529_),
    .ZN(_2758_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _7625_ (.A1(_2756_),
    .A2(_2749_),
    .B(_2758_),
    .ZN(_2759_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _7626_ (.A1(_0933_),
    .A2(_0594_),
    .Z(_2760_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _7627_ (.A1(_2760_),
    .A2(_2697_),
    .B(_2728_),
    .ZN(_2761_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _7628_ (.A1(_2727_),
    .A2(_2761_),
    .ZN(_2762_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7629_ (.A1(_1680_),
    .A2(_2762_),
    .ZN(_2763_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7630_ (.A1(_2757_),
    .A2(_1614_),
    .ZN(_2764_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _7631_ (.A1(_2499_),
    .A2(_2763_),
    .A3(_2764_),
    .ZN(_2765_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7632_ (.A1(_2759_),
    .A2(_2765_),
    .ZN(_2766_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _7633_ (.A1(_0940_),
    .A2(_2655_),
    .B1(_2766_),
    .B2(_1443_),
    .ZN(_2767_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _7634_ (.A1(_2196_),
    .A2(_2686_),
    .B1(_2753_),
    .B2(_2767_),
    .ZN(_2768_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _7635_ (.A1(_2752_),
    .A2(_2768_),
    .B(_2573_),
    .ZN(_2769_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _7636_ (.A1(_2197_),
    .A2(_2580_),
    .B(_2769_),
    .ZN(_2770_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7637_ (.I(_2465_),
    .Z(_2771_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7638_ (.I(_1634_),
    .Z(_2772_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _7639_ (.A1(_2757_),
    .A2(_2771_),
    .B(_2772_),
    .ZN(_2773_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _7640_ (.A1(_2579_),
    .A2(_2770_),
    .B(_2773_),
    .ZN(_0178_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7641_ (.I(_2520_),
    .Z(_2774_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7642_ (.A1(_0948_),
    .A2(_2655_),
    .ZN(_2775_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7643_ (.I(_2503_),
    .Z(_2776_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _7644_ (.I(_2776_),
    .Z(_2777_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _7645_ (.I(net34),
    .Z(_2778_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7646_ (.A1(_2757_),
    .A2(_2747_),
    .ZN(_2779_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _7647_ (.A1(_2778_),
    .A2(_2779_),
    .Z(_2780_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_1 _7648_ (.A1(_2778_),
    .A2(_2531_),
    .B1(_2534_),
    .B2(_1526_),
    .C(_2501_),
    .ZN(_2781_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _7649_ (.A1(_2777_),
    .A2(_2780_),
    .B(_2781_),
    .ZN(_2782_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _7650_ (.A1(\as2650.pc[6] ),
    .A2(net2),
    .Z(_2783_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _7651_ (.I(_2783_),
    .ZN(_2784_));
 gf180mcu_fd_sc_mcu7t5v0__or4_1 _7652_ (.A1(_2636_),
    .A2(_2760_),
    .A3(_2696_),
    .A4(_2726_),
    .Z(_2785_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7653_ (.A1(_2194_),
    .A2(_0682_),
    .ZN(_2786_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _7654_ (.A1(_2194_),
    .A2(net1),
    .B(net10),
    .C(_2187_),
    .ZN(_2787_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _7655_ (.A1(_2786_),
    .A2(_2787_),
    .Z(_2788_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7656_ (.A1(_2785_),
    .A2(_2788_),
    .ZN(_2789_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _7657_ (.A1(_2784_),
    .A2(_2789_),
    .Z(_2790_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _7658_ (.A1(_2778_),
    .A2(_2542_),
    .B(_2499_),
    .ZN(_2791_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _7659_ (.A1(_1619_),
    .A2(_2790_),
    .B(_2791_),
    .ZN(_2792_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7660_ (.I(_1271_),
    .Z(_2793_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7661_ (.I(_2793_),
    .Z(_2794_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _7662_ (.A1(_2782_),
    .A2(_2792_),
    .B(_2794_),
    .ZN(_2795_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7663_ (.A1(_2632_),
    .A2(_2795_),
    .ZN(_2796_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _7664_ (.A1(_0948_),
    .A2(_2686_),
    .B(_2796_),
    .ZN(_2797_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _7665_ (.A1(_1587_),
    .A2(_0748_),
    .Z(_2798_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _7666_ (.A1(_0682_),
    .A2(_0667_),
    .Z(_2799_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7667_ (.I(_0682_),
    .Z(_2800_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _7668_ (.A1(_2800_),
    .A2(_0667_),
    .Z(_2801_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _7669_ (.A1(_2799_),
    .A2(_2734_),
    .B(_2801_),
    .ZN(_2802_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _7670_ (.A1(_2798_),
    .A2(_2802_),
    .ZN(_2803_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7671_ (.A1(_2555_),
    .A2(_2803_),
    .ZN(_2804_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _7672_ (.A1(_1559_),
    .A2(_2553_),
    .B(_2467_),
    .C(_2804_),
    .ZN(_2805_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _7673_ (.A1(_1587_),
    .A2(_0770_),
    .Z(_2806_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _7674_ (.A1(_2800_),
    .A2(_0697_),
    .Z(_2807_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _7675_ (.A1(_0683_),
    .A2(_0697_),
    .Z(_2808_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _7676_ (.A1(_2807_),
    .A2(_2741_),
    .B(_2808_),
    .ZN(_2809_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _7677_ (.A1(_2806_),
    .A2(_2809_),
    .ZN(_2810_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7678_ (.A1(_2473_),
    .A2(_2810_),
    .ZN(_2811_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _7679_ (.A1(_1559_),
    .A2(_2560_),
    .B(_2811_),
    .C(_2565_),
    .ZN(_2812_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _7680_ (.A1(_2805_),
    .A2(_2812_),
    .B(_1311_),
    .ZN(_2813_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7681_ (.A1(_2786_),
    .A2(_2787_),
    .ZN(_2814_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _7682_ (.A1(_2729_),
    .A2(_2727_),
    .ZN(_2815_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _7683_ (.A1(_2814_),
    .A2(_2815_),
    .ZN(_2816_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _7684_ (.A1(_2783_),
    .A2(_2816_),
    .Z(_2817_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7685_ (.I(_2485_),
    .Z(_2818_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _7686_ (.A1(_2613_),
    .A2(_2780_),
    .B1(_2817_),
    .B2(_2818_),
    .ZN(_2819_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _7687_ (.A1(_2751_),
    .A2(_2813_),
    .A3(_2819_),
    .ZN(_2820_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _7688_ (.A1(_2775_),
    .A2(_2797_),
    .B(_2820_),
    .ZN(_2821_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _7689_ (.A1(_2201_),
    .A2(_2684_),
    .B1(_2821_),
    .B2(_2681_),
    .ZN(_2822_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _7690_ (.A1(_2778_),
    .A2(_2771_),
    .B(_2772_),
    .ZN(_2823_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _7691_ (.A1(_2774_),
    .A2(_2822_),
    .B(_2823_),
    .ZN(_0179_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _7692_ (.I(_2573_),
    .Z(_2824_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _7693_ (.I(_0756_),
    .Z(_2825_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7694_ (.A1(_2825_),
    .A2(_0749_),
    .ZN(_2826_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _7695_ (.A1(_2798_),
    .A2(_2802_),
    .B(_2826_),
    .ZN(_2827_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _7696_ (.A1(_1617_),
    .A2(_0828_),
    .A3(_2827_),
    .Z(_2828_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7697_ (.A1(_1680_),
    .A2(_2588_),
    .ZN(_2829_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _7698_ (.A1(_2588_),
    .A2(_2828_),
    .B(_2829_),
    .C(_2554_),
    .ZN(_2830_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7699_ (.A1(_0757_),
    .A2(_0771_),
    .ZN(_2831_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _7700_ (.A1(_2806_),
    .A2(_2809_),
    .B(_2831_),
    .ZN(_2832_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _7701_ (.A1(_1599_),
    .A2(_0830_),
    .A3(_2832_),
    .Z(_2833_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7702_ (.A1(_1680_),
    .A2(_2704_),
    .ZN(_2834_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _7703_ (.A1(_2704_),
    .A2(_2833_),
    .B(_2834_),
    .C(_2476_),
    .ZN(_2835_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _7704_ (.I(_1330_),
    .Z(_2836_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _7705_ (.A1(_2830_),
    .A2(_2835_),
    .B(_2836_),
    .ZN(_2837_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _7706_ (.I(net54),
    .ZN(_2838_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _7707_ (.A1(net34),
    .A2(net33),
    .A3(_2747_),
    .ZN(_2839_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _7708_ (.A1(_2838_),
    .A2(_2839_),
    .Z(_2840_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _7709_ (.A1(_2720_),
    .A2(_2840_),
    .B(_2818_),
    .ZN(_2841_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _7710_ (.A1(\as2650.pc[7] ),
    .A2(net2),
    .Z(_2842_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7711_ (.A1(_0945_),
    .A2(net2),
    .ZN(_2843_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _7712_ (.A1(_2784_),
    .A2(_2816_),
    .B(_2843_),
    .ZN(_2844_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _7713_ (.A1(_2842_),
    .A2(_2844_),
    .ZN(_2845_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _7714_ (.A1(_2837_),
    .A2(_2841_),
    .B1(_2845_),
    .B2(_2818_),
    .ZN(_2846_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7715_ (.A1(_2783_),
    .A2(_2789_),
    .ZN(_2847_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7716_ (.A1(_2843_),
    .A2(_2847_),
    .ZN(_2848_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _7717_ (.A1(_2842_),
    .A2(_2848_),
    .Z(_2849_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7718_ (.A1(_2618_),
    .A2(_2849_),
    .ZN(_2850_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _7719_ (.A1(_2491_),
    .A2(_2646_),
    .ZN(_2851_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7720_ (.A1(_1516_),
    .A2(_2851_),
    .ZN(_2852_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _7721_ (.A1(net54),
    .A2(_2644_),
    .B(_2852_),
    .ZN(_2853_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7722_ (.I(_1479_),
    .Z(_2854_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _7723_ (.A1(_1497_),
    .A2(_1683_),
    .ZN(_2855_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7724_ (.I(_2855_),
    .Z(_2856_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7725_ (.A1(_2648_),
    .A2(_2840_),
    .ZN(_2857_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _7726_ (.A1(net54),
    .A2(_2505_),
    .B1(_2688_),
    .B2(_2542_),
    .ZN(_2858_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _7727_ (.A1(_2854_),
    .A2(_2856_),
    .A3(_2857_),
    .A4(_2858_),
    .ZN(_2859_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _7728_ (.A1(_2204_),
    .A2(_2496_),
    .B(_2859_),
    .ZN(_2860_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _7729_ (.A1(_2850_),
    .A2(_2853_),
    .B1(_2860_),
    .B2(_1450_),
    .ZN(_2861_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _7730_ (.A1(_2751_),
    .A2(_2846_),
    .B(_2861_),
    .ZN(_2862_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7731_ (.A1(_2824_),
    .A2(_2862_),
    .ZN(_2863_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _7732_ (.A1(_2205_),
    .A2(_2580_),
    .B(_2863_),
    .ZN(_2864_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _7733_ (.A1(net54),
    .A2(_2771_),
    .B(_2772_),
    .ZN(_2865_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _7734_ (.A1(_2774_),
    .A2(_2864_),
    .B(_2865_),
    .ZN(_0180_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7735_ (.I(\as2650.addr_buff[0] ),
    .Z(_2866_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_2 _7736_ (.A1(_0835_),
    .A2(_0827_),
    .B1(_2798_),
    .B2(_2802_),
    .C(_2826_),
    .ZN(_2867_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _7737_ (.A1(_0836_),
    .A2(_0827_),
    .B(_4245_),
    .ZN(_2868_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7738_ (.I(_2868_),
    .Z(_2869_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _7739_ (.A1(_2866_),
    .A2(_2867_),
    .A3(_2869_),
    .ZN(_2870_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7740_ (.I(_2867_),
    .Z(_2871_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7741_ (.A1(_2871_),
    .A2(_2869_),
    .ZN(_2872_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7742_ (.A1(_2334_),
    .A2(_2872_),
    .ZN(_2873_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7743_ (.A1(_2870_),
    .A2(_2873_),
    .ZN(_2874_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7744_ (.A1(_1616_),
    .A2(_0829_),
    .ZN(_2875_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_2 _7745_ (.A1(_2806_),
    .A2(_2809_),
    .B(_2875_),
    .C(_2831_),
    .ZN(_2876_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _7746_ (.A1(_1604_),
    .A2(_0829_),
    .ZN(_2877_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _7747_ (.A1(_2703_),
    .A2(_2877_),
    .ZN(_2878_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _7748_ (.A1(_2866_),
    .A2(_2876_),
    .A3(_2878_),
    .ZN(_2879_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7749_ (.A1(_2876_),
    .A2(_2878_),
    .ZN(_2880_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7750_ (.A1(_2334_),
    .A2(_2880_),
    .ZN(_2881_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7751_ (.A1(_2879_),
    .A2(_2881_),
    .ZN(_2882_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _7752_ (.A1(_2467_),
    .A2(_2874_),
    .B1(_2882_),
    .B2(_2598_),
    .ZN(_2883_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _7753_ (.I(net36),
    .Z(_2884_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _7754_ (.A1(_2838_),
    .A2(_2839_),
    .ZN(_2885_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _7755_ (.A1(_2884_),
    .A2(_2885_),
    .ZN(_2886_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7756_ (.A1(_2480_),
    .A2(_2886_),
    .ZN(_2887_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _7757_ (.I(_2485_),
    .Z(_2888_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _7758_ (.A1(_2836_),
    .A2(_2883_),
    .B(_2887_),
    .C(_2888_),
    .ZN(_2889_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _7759_ (.A1(\as2650.pc[8] ),
    .A2(_0755_),
    .Z(_2890_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7760_ (.A1(_2783_),
    .A2(_2842_),
    .ZN(_2891_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _7761_ (.A1(_2788_),
    .A2(_2891_),
    .B(_2843_),
    .ZN(_2892_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _7762_ (.A1(_2203_),
    .A2(_0755_),
    .B(_2892_),
    .ZN(_2893_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_1 _7763_ (.A1(_2729_),
    .A2(_2727_),
    .A3(_2891_),
    .B(_2893_),
    .ZN(_2894_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7764_ (.A1(_2890_),
    .A2(_2894_),
    .ZN(_2895_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _7765_ (.A1(_2890_),
    .A2(_2894_),
    .B(_2607_),
    .ZN(_2896_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _7766_ (.I(_2896_),
    .ZN(_2897_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _7767_ (.A1(_2895_),
    .A2(_2897_),
    .B(_2751_),
    .ZN(_2898_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _7768_ (.I(_2866_),
    .Z(_2899_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_1 _7769_ (.A1(_2884_),
    .A2(_2532_),
    .B1(_2535_),
    .B2(_2899_),
    .C(_2502_),
    .ZN(_2900_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _7770_ (.A1(_2386_),
    .A2(_2886_),
    .B(_2900_),
    .ZN(_2901_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _7771_ (.A1(_2785_),
    .A2(_2891_),
    .B(_2893_),
    .ZN(_2902_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _7772_ (.A1(_2890_),
    .A2(_2902_),
    .ZN(_2903_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _7773_ (.A1(_2884_),
    .A2(_2618_),
    .B(_2500_),
    .ZN(_2904_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _7774_ (.A1(_1546_),
    .A2(_2903_),
    .B(_2904_),
    .ZN(_2905_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _7775_ (.A1(_2901_),
    .A2(_2905_),
    .B(_2550_),
    .ZN(_2906_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _7776_ (.A1(_0966_),
    .A2(_2528_),
    .B(_2624_),
    .ZN(_2907_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _7777_ (.A1(_2889_),
    .A2(_2898_),
    .B1(_2906_),
    .B2(_2907_),
    .ZN(_2908_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _7778_ (.A1(_0966_),
    .A2(_2684_),
    .B1(_2908_),
    .B2(_2681_),
    .ZN(_2909_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _7779_ (.A1(_2884_),
    .A2(_2771_),
    .B(_2772_),
    .ZN(_2910_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _7780_ (.A1(_2774_),
    .A2(_2909_),
    .B(_2910_),
    .ZN(_0181_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _7781_ (.I(\as2650.pc[9] ),
    .ZN(_2911_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _7782_ (.A1(_2911_),
    .A2(_1586_),
    .Z(_2912_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7783_ (.A1(_0964_),
    .A2(_0757_),
    .ZN(_2913_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7784_ (.A1(_2913_),
    .A2(_2895_),
    .ZN(_2914_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _7785_ (.A1(_2912_),
    .A2(_2914_),
    .Z(_2915_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _7786_ (.A1(_2361_),
    .A2(_2879_),
    .Z(_2916_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _7787_ (.A1(_2361_),
    .A2(_2870_),
    .Z(_2917_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _7788_ (.A1(_2476_),
    .A2(_2916_),
    .B1(_2917_),
    .B2(_2554_),
    .ZN(_2918_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _7789_ (.I(net37),
    .Z(_2919_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7790_ (.A1(net36),
    .A2(_2885_),
    .ZN(_2920_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _7791_ (.A1(_2919_),
    .A2(_2920_),
    .ZN(_2921_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_1 _7792_ (.A1(_2836_),
    .A2(_2918_),
    .B1(_2921_),
    .B2(_2720_),
    .C(_2486_),
    .ZN(_2922_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7793_ (.I(_2570_),
    .Z(_2923_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _7794_ (.A1(_2818_),
    .A2(_2915_),
    .B(_2922_),
    .C(_2923_),
    .ZN(_2924_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7795_ (.I(_1479_),
    .Z(_2925_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7796_ (.I(_2925_),
    .Z(_2926_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7797_ (.I(_2855_),
    .Z(_2927_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7798_ (.I(_2927_),
    .Z(_2928_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7799_ (.A1(_2777_),
    .A2(_2921_),
    .ZN(_2929_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _7800_ (.A1(_2919_),
    .A2(_2505_),
    .B1(_2688_),
    .B2(_2362_),
    .ZN(_2930_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _7801_ (.A1(_2926_),
    .A2(_2928_),
    .A3(_2929_),
    .A4(_2930_),
    .ZN(_2931_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _7802_ (.A1(_0979_),
    .A2(_2496_),
    .B(_2931_),
    .ZN(_2932_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7803_ (.A1(_2514_),
    .A2(_2932_),
    .ZN(_2933_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7804_ (.A1(_2890_),
    .A2(_2902_),
    .ZN(_2934_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7805_ (.A1(_2913_),
    .A2(_2934_),
    .ZN(_2935_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _7806_ (.A1(_2912_),
    .A2(_2935_),
    .Z(_2936_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _7807_ (.A1(_2919_),
    .A2(_2644_),
    .B(_2852_),
    .ZN(_2937_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _7808_ (.A1(_2377_),
    .A2(_2936_),
    .B(_2937_),
    .ZN(_2938_));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _7809_ (.A1(_2924_),
    .A2(_2933_),
    .A3(_2938_),
    .Z(_2939_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7810_ (.I(_1327_),
    .Z(_2940_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _7811_ (.A1(_0979_),
    .A2(_2684_),
    .B1(_2939_),
    .B2(_2940_),
    .ZN(_2941_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7812_ (.I(_2465_),
    .Z(_2942_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7813_ (.I(_1565_),
    .Z(_2943_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _7814_ (.A1(_2919_),
    .A2(_2942_),
    .B(_2943_),
    .ZN(_2944_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _7815_ (.A1(_2774_),
    .A2(_2941_),
    .B(_2944_),
    .ZN(_0182_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _7816_ (.I(net53),
    .ZN(_2945_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _7817_ (.A1(net37),
    .A2(net36),
    .A3(_2885_),
    .ZN(_2946_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _7818_ (.A1(_2945_),
    .A2(_2946_),
    .Z(_2947_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _7819_ (.A1(_2744_),
    .A2(_2876_),
    .A3(_2878_),
    .ZN(_2948_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _7820_ (.A1(_2662_),
    .A2(_2871_),
    .A3(_2869_),
    .ZN(_2949_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _7821_ (.A1(_2899_),
    .A2(_2361_),
    .A3(_2366_),
    .ZN(_2950_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _7822_ (.A1(_2948_),
    .A2(_2949_),
    .B(_2950_),
    .ZN(_2951_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7823_ (.A1(_2866_),
    .A2(\as2650.addr_buff[1] ),
    .ZN(_2952_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _7824_ (.A1(_2871_),
    .A2(_2869_),
    .B(_2564_),
    .ZN(_2953_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _7825_ (.A1(_2336_),
    .A2(_2612_),
    .B1(_2952_),
    .B2(_2953_),
    .ZN(_2954_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _7826_ (.A1(_2880_),
    .A2(_2952_),
    .B(_2744_),
    .ZN(_2955_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _7827_ (.A1(_2954_),
    .A2(_2955_),
    .B(_2366_),
    .ZN(_2956_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _7828_ (.A1(_2951_),
    .A2(_2956_),
    .B(_2661_),
    .ZN(_2957_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _7829_ (.A1(_2613_),
    .A2(_2947_),
    .B(_2957_),
    .C(_2888_),
    .ZN(_2958_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _7830_ (.A1(\as2650.pc[10] ),
    .A2(_1586_),
    .Z(_2959_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7831_ (.I(_2959_),
    .Z(_2960_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _7832_ (.A1(\as2650.pc[9] ),
    .A2(_0964_),
    .B(_0756_),
    .ZN(_2961_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _7833_ (.I(_2961_),
    .ZN(_2962_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _7834_ (.A1(_2895_),
    .A2(_2912_),
    .ZN(_2963_));
 gf180mcu_fd_sc_mcu7t5v0__or3_1 _7835_ (.A1(_2960_),
    .A2(_2962_),
    .A3(_2963_),
    .Z(_2964_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _7836_ (.A1(_2962_),
    .A2(_2963_),
    .B(_2960_),
    .ZN(_2965_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _7837_ (.A1(_2658_),
    .A2(_2964_),
    .A3(_2965_),
    .ZN(_2966_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _7838_ (.A1(_2923_),
    .A2(_2966_),
    .Z(_2967_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _7839_ (.I(_0988_),
    .ZN(_2968_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _7840_ (.I(_2968_),
    .Z(_2969_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _7841_ (.A1(_2540_),
    .A2(_2947_),
    .ZN(_2970_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_1 _7842_ (.A1(net53),
    .A2(_2531_),
    .B1(_2535_),
    .B2(_2366_),
    .C(_2854_),
    .ZN(_2971_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _7843_ (.A1(_2969_),
    .A2(_2527_),
    .B1(_2970_),
    .B2(_2971_),
    .ZN(_2972_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _7844_ (.A1(_0990_),
    .A2(_2513_),
    .B1(_2972_),
    .B2(_2928_),
    .C(_2551_),
    .ZN(_2973_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _7845_ (.A1(_2934_),
    .A2(_2912_),
    .Z(_2974_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7846_ (.A1(_2961_),
    .A2(_2974_),
    .ZN(_2975_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _7847_ (.A1(_2960_),
    .A2(_2975_),
    .ZN(_2976_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7848_ (.A1(_1546_),
    .A2(_2976_),
    .ZN(_2977_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _7849_ (.A1(net53),
    .A2(_1711_),
    .B(_2851_),
    .C(_2977_),
    .ZN(_2978_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _7850_ (.A1(_2958_),
    .A2(_2967_),
    .B1(_2973_),
    .B2(_2978_),
    .ZN(_2979_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _7851_ (.A1(_0990_),
    .A2(_2522_),
    .B1(_2979_),
    .B2(_2940_),
    .ZN(_2980_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _7852_ (.A1(net53),
    .A2(_2942_),
    .B(_2943_),
    .ZN(_2981_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _7853_ (.A1(_2521_),
    .A2(_2980_),
    .B(_2981_),
    .ZN(_0183_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7854_ (.I(net39),
    .Z(_2982_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _7855_ (.A1(_2945_),
    .A2(_2946_),
    .ZN(_2983_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _7856_ (.A1(_2982_),
    .A2(_2983_),
    .Z(_2984_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _7857_ (.A1(_2953_),
    .A2(_2950_),
    .B(_2612_),
    .ZN(_2985_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _7858_ (.A1(_2880_),
    .A2(_2950_),
    .B(_2744_),
    .ZN(_2986_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _7859_ (.A1(_2369_),
    .A2(_2985_),
    .A3(_2986_),
    .ZN(_2987_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _7860_ (.A1(_2369_),
    .A2(_2951_),
    .B(_2987_),
    .C(_2661_),
    .ZN(_2988_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _7861_ (.A1(_2613_),
    .A2(_2984_),
    .B(_2988_),
    .C(_2888_),
    .ZN(_2989_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _7862_ (.A1(\as2650.pc[11] ),
    .A2(_1586_),
    .Z(_2990_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7863_ (.A1(_0989_),
    .A2(_0757_),
    .ZN(_2991_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7864_ (.A1(_2991_),
    .A2(_2965_),
    .ZN(_2992_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _7865_ (.A1(_2990_),
    .A2(_2992_),
    .Z(_2993_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _7866_ (.A1(_2719_),
    .A2(_2993_),
    .B(_2483_),
    .ZN(_2994_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _7867_ (.I(_0997_),
    .ZN(_2995_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7868_ (.I(_2494_),
    .Z(_2996_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7869_ (.A1(_2385_),
    .A2(_2984_),
    .ZN(_2997_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _7870_ (.I(\as2650.addr_buff[3] ),
    .Z(_2998_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _7871_ (.A1(_2982_),
    .A2(_2504_),
    .B1(_2507_),
    .B2(_2998_),
    .C(_1268_),
    .ZN(_2999_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _7872_ (.A1(_2995_),
    .A2(_2996_),
    .B1(_2997_),
    .B2(_2999_),
    .ZN(_3000_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7873_ (.I(_2149_),
    .Z(_3001_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _7874_ (.A1(_0997_),
    .A2(_2525_),
    .B1(_3000_),
    .B2(_3001_),
    .ZN(_3002_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _7875_ (.A1(_1575_),
    .A2(_3002_),
    .Z(_3003_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7876_ (.A1(_2960_),
    .A2(_2975_),
    .ZN(_3004_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7877_ (.A1(_2991_),
    .A2(_3004_),
    .ZN(_3005_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _7878_ (.A1(_2990_),
    .A2(_3005_),
    .Z(_3006_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _7879_ (.A1(_2982_),
    .A2(_2644_),
    .Z(_3007_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _7880_ (.A1(_1546_),
    .A2(_3006_),
    .B(_3007_),
    .C(_2852_),
    .ZN(_3008_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _7881_ (.A1(_2989_),
    .A2(_2994_),
    .B(_3003_),
    .C(_3008_),
    .ZN(_3009_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _7882_ (.A1(_0997_),
    .A2(_2522_),
    .B1(_3009_),
    .B2(_2940_),
    .ZN(_3010_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _7883_ (.A1(_2982_),
    .A2(_2942_),
    .B(_2943_),
    .ZN(_3011_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _7884_ (.A1(_2521_),
    .A2(_3010_),
    .B(_3011_),
    .ZN(_0184_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _7885_ (.A1(\as2650.pc[12] ),
    .A2(_0756_),
    .Z(_3012_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _7886_ (.A1(_2959_),
    .A2(_2990_),
    .Z(_3013_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _7887_ (.I(_3013_),
    .ZN(_3014_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _7888_ (.A1(\as2650.pc[11] ),
    .A2(_0988_),
    .B(_2825_),
    .ZN(_3015_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _7889_ (.A1(_2974_),
    .A2(_3014_),
    .B(_3015_),
    .C(_2961_),
    .ZN(_3016_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _7890_ (.A1(_3012_),
    .A2(_3016_),
    .Z(_3017_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7891_ (.A1(_1711_),
    .A2(_3017_),
    .ZN(_3018_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _7892_ (.A1(net52),
    .A2(_2377_),
    .B(_2852_),
    .ZN(_3019_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _7893_ (.I(\as2650.addr_buff[4] ),
    .Z(_3020_));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _7894_ (.A1(\as2650.addr_buff[0] ),
    .A2(\as2650.addr_buff[1] ),
    .A3(\as2650.addr_buff[2] ),
    .Z(_3021_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _7895_ (.A1(_2998_),
    .A2(_2871_),
    .A3(_2868_),
    .A4(_3021_),
    .ZN(_3022_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _7896_ (.A1(_3020_),
    .A2(_3022_),
    .Z(_3023_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _7897_ (.A1(_2998_),
    .A2(_2876_),
    .A3(_2878_),
    .A4(_3021_),
    .ZN(_3024_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _7898_ (.A1(_3020_),
    .A2(_3024_),
    .Z(_3025_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _7899_ (.A1(_2662_),
    .A2(_3023_),
    .B1(_3025_),
    .B2(_2476_),
    .ZN(_3026_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7900_ (.A1(net39),
    .A2(_2983_),
    .ZN(_3027_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _7901_ (.A1(net52),
    .A2(_3027_),
    .ZN(_3028_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_1 _7902_ (.A1(_2836_),
    .A2(_3026_),
    .B1(_3028_),
    .B2(_2720_),
    .C(_2486_),
    .ZN(_3029_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7903_ (.A1(_2961_),
    .A2(_3015_),
    .ZN(_3030_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _7904_ (.A1(_2963_),
    .A2(_3013_),
    .B(_3030_),
    .ZN(_3031_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _7905_ (.A1(_3012_),
    .A2(_3031_),
    .ZN(_3032_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7906_ (.A1(_2607_),
    .A2(_3032_),
    .ZN(_3033_));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _7907_ (.A1(_2923_),
    .A2(_3029_),
    .A3(_3033_),
    .Z(_3034_));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _7908_ (.I(\as2650.pc[12] ),
    .ZN(_3035_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7909_ (.A1(_2385_),
    .A2(_3028_),
    .ZN(_3036_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _7910_ (.A1(net52),
    .A2(_2504_),
    .B1(_2507_),
    .B2(_3020_),
    .C(_1268_),
    .ZN(_3037_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _7911_ (.A1(_3035_),
    .A2(_2495_),
    .B1(_3036_),
    .B2(_3037_),
    .ZN(_3038_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _7912_ (.A1(_1003_),
    .A2(_2525_),
    .B1(_3038_),
    .B2(_3001_),
    .ZN(_3039_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _7913_ (.A1(_1450_),
    .A2(_3039_),
    .Z(_3040_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _7914_ (.A1(_3018_),
    .A2(_3019_),
    .B(_3034_),
    .C(_3040_),
    .ZN(_3041_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _7915_ (.A1(_1003_),
    .A2(_2522_),
    .B1(_3041_),
    .B2(_2940_),
    .ZN(_3042_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _7916_ (.A1(net52),
    .A2(_2942_),
    .B(_2943_),
    .ZN(_3043_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _7917_ (.A1(_2521_),
    .A2(_3042_),
    .B(_3043_),
    .ZN(_0185_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _7918_ (.I(_2445_),
    .ZN(_3044_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7919_ (.I(_1320_),
    .Z(_3045_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _7920_ (.A1(_1462_),
    .A2(_1327_),
    .ZN(_3046_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _7921_ (.A1(_3045_),
    .A2(_2354_),
    .A3(_3046_),
    .A4(_2433_),
    .ZN(_3047_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7922_ (.I(_0871_),
    .Z(_3048_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _7923_ (.A1(_3048_),
    .A2(_2152_),
    .B(_4444_),
    .ZN(_3049_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_2 _7924_ (.A1(_1331_),
    .A2(_2412_),
    .A3(_3047_),
    .A4(_3049_),
    .ZN(_3050_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7925_ (.A1(_1480_),
    .A2(_2427_),
    .ZN(_3051_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _7926_ (.A1(_2457_),
    .A2(_2425_),
    .A3(_3051_),
    .ZN(_3052_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7927_ (.A1(_4491_),
    .A2(_2446_),
    .ZN(_3053_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_2 _7928_ (.A1(_1353_),
    .A2(_3050_),
    .A3(_3052_),
    .A4(_3053_),
    .ZN(_3054_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _7929_ (.A1(_2422_),
    .A2(_2453_),
    .Z(_3055_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_2 _7930_ (.A1(_3044_),
    .A2(_2462_),
    .A3(_3054_),
    .A4(_3055_),
    .ZN(_3056_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7931_ (.I(_2157_),
    .Z(_3057_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7932_ (.I(_3057_),
    .Z(_3058_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _7933_ (.I(_3058_),
    .Z(_3059_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _7934_ (.A1(_2551_),
    .A2(_4187_),
    .A3(_3059_),
    .ZN(_3060_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7935_ (.I(_1324_),
    .Z(_3061_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_1 _7936_ (.A1(net26),
    .A2(_1367_),
    .B1(_3061_),
    .B2(_1575_),
    .C(_1443_),
    .ZN(_3062_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _7937_ (.A1(_2686_),
    .A2(_2381_),
    .B1(_3060_),
    .B2(_3062_),
    .ZN(_3063_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _7938_ (.A1(_2824_),
    .A2(_3063_),
    .B(_3056_),
    .ZN(_3064_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _7939_ (.A1(net49),
    .A2(_3056_),
    .B(_3064_),
    .C(_2578_),
    .ZN(_0186_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_2 _7940_ (.A1(_1356_),
    .A2(_1684_),
    .A3(_1504_),
    .ZN(_3065_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _7941_ (.A1(_4169_),
    .A2(_2348_),
    .ZN(_3066_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _7942_ (.A1(_0891_),
    .A2(_3066_),
    .ZN(_3067_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7943_ (.A1(_3065_),
    .A2(_3067_),
    .ZN(_3068_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _7944_ (.A1(_2349_),
    .A2(_3068_),
    .ZN(_3069_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _7945_ (.I(_2347_),
    .Z(_3070_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_2 _7946_ (.A1(_4237_),
    .A2(_2348_),
    .A3(_3070_),
    .ZN(_3071_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _7947_ (.A1(_3069_),
    .A2(_3071_),
    .ZN(_3072_));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _7948_ (.A1(_4490_),
    .A2(_2444_),
    .A3(_2446_),
    .Z(_3073_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _7949_ (.I(_1503_),
    .Z(_3074_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _7950_ (.A1(_2450_),
    .A2(_3074_),
    .A3(_2412_),
    .A4(_2451_),
    .ZN(_3075_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7951_ (.I(_2157_),
    .Z(_3076_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _7952_ (.A1(_2396_),
    .A2(_3076_),
    .B1(_2407_),
    .B2(_1163_),
    .C(_1319_),
    .ZN(_3077_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _7953_ (.A1(_1087_),
    .A2(_2441_),
    .A3(_3077_),
    .ZN(_3078_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _7954_ (.A1(_2426_),
    .A2(_3075_),
    .A3(_3078_),
    .ZN(_3079_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _7955_ (.I(_1516_),
    .Z(_3080_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7956_ (.A1(_1617_),
    .A2(_2352_),
    .ZN(_3081_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _7957_ (.I(_2493_),
    .Z(_3082_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _7958_ (.A1(_1482_),
    .A2(_1293_),
    .A3(_2160_),
    .A4(_3082_),
    .ZN(_3083_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _7959_ (.A1(_2149_),
    .A2(_3081_),
    .B(_3083_),
    .ZN(_3084_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7960_ (.A1(_3080_),
    .A2(_3084_),
    .ZN(_3085_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _7961_ (.A1(_3072_),
    .A2(_3073_),
    .A3(_3079_),
    .A4(_3085_),
    .ZN(_3086_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _7962_ (.A1(_2463_),
    .A2(_3086_),
    .ZN(_3087_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _7963_ (.I(_1517_),
    .Z(_3088_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _7964_ (.I(_1275_),
    .Z(_3089_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7965_ (.I(_3089_),
    .Z(_3090_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7966_ (.A1(net51),
    .A2(_3090_),
    .ZN(_3091_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _7967_ (.A1(_2380_),
    .A2(_3091_),
    .B(_1481_),
    .ZN(_3092_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7968_ (.I(_2160_),
    .Z(_3093_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _7969_ (.A1(_3093_),
    .A2(_2155_),
    .B(_2508_),
    .ZN(_3094_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7970_ (.I(_0872_),
    .Z(_3095_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _7971_ (.A1(net51),
    .A2(_1277_),
    .A3(_3095_),
    .ZN(_3096_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _7972_ (.A1(_3094_),
    .A2(_3096_),
    .B(_1686_),
    .C(_2525_),
    .ZN(_3097_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7973_ (.A1(_3092_),
    .A2(_3097_),
    .ZN(_3098_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _7974_ (.A1(net51),
    .A2(_3090_),
    .A3(_2155_),
    .ZN(_3099_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _7975_ (.A1(_3088_),
    .A2(_3098_),
    .B1(_3099_),
    .B2(_2923_),
    .ZN(_3100_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _7976_ (.A1(_1692_),
    .A2(_3100_),
    .B(_2403_),
    .ZN(_3101_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _7977_ (.A1(net51),
    .A2(_3087_),
    .ZN(_3102_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _7978_ (.A1(_3087_),
    .A2(_3101_),
    .B(_3102_),
    .C(_2578_),
    .ZN(_0187_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _7979_ (.I(_2793_),
    .Z(_3103_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _7980_ (.A1(_3103_),
    .A2(_2338_),
    .A3(_1312_),
    .ZN(_3104_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7981_ (.A1(_2551_),
    .A2(_3104_),
    .ZN(_3105_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _7982_ (.I(_1486_),
    .Z(_3106_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_4 _7983_ (.A1(_2407_),
    .A2(_3105_),
    .B(_2434_),
    .C(_3106_),
    .ZN(_3107_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7984_ (.A1(_4265_),
    .A2(_2824_),
    .ZN(_3108_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _7985_ (.A1(_4244_),
    .A2(_3107_),
    .ZN(_3109_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _7986_ (.A1(_3107_),
    .A2(_3108_),
    .B(_3109_),
    .C(_2578_),
    .ZN(_0188_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7987_ (.A1(_4264_),
    .A2(_2824_),
    .ZN(_3110_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _7988_ (.A1(_4243_),
    .A2(_3107_),
    .ZN(_3111_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _7989_ (.I(_2577_),
    .Z(_3112_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _7990_ (.A1(_3107_),
    .A2(_3110_),
    .B(_3111_),
    .C(_3112_),
    .ZN(_0189_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7991_ (.A1(_4406_),
    .A2(_1524_),
    .ZN(_3113_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7992_ (.A1(_1550_),
    .A2(_1442_),
    .ZN(_3114_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7993_ (.A1(_3113_),
    .A2(_3114_),
    .ZN(_3115_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7994_ (.A1(_1367_),
    .A2(_2420_),
    .ZN(_3116_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _7995_ (.A1(_1457_),
    .A2(_1477_),
    .B(_1571_),
    .ZN(_3117_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_2 _7996_ (.A1(_1277_),
    .A2(_1493_),
    .B(_1517_),
    .C(_0852_),
    .ZN(_3118_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _7997_ (.A1(_3116_),
    .A2(_3117_),
    .A3(_3118_),
    .ZN(_3119_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _7998_ (.I(_3119_),
    .Z(_3120_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _7999_ (.I0(_3115_),
    .I1(_4291_),
    .S(_3120_),
    .Z(_3121_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _8000_ (.I(_3121_),
    .Z(_0190_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _8001_ (.A1(_2536_),
    .A2(_1289_),
    .ZN(_3122_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _8002_ (.A1(_4542_),
    .A2(_1294_),
    .ZN(_3123_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _8003_ (.A1(_3122_),
    .A2(_3123_),
    .ZN(_3124_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _8004_ (.I0(_3124_),
    .I1(_0297_),
    .S(_3120_),
    .Z(_3125_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _8005_ (.I(_3125_),
    .Z(_0191_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _8006_ (.I(_1289_),
    .Z(_3126_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _8007_ (.A1(_0361_),
    .A2(_3126_),
    .ZN(_3127_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _8008_ (.A1(_1699_),
    .A2(_1295_),
    .ZN(_3128_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _8009_ (.A1(_3127_),
    .A2(_3128_),
    .ZN(_3129_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _8010_ (.I(_3119_),
    .Z(_3130_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _8011_ (.I0(_3129_),
    .I1(_0413_),
    .S(_3130_),
    .Z(_3131_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _8012_ (.I(_3131_),
    .Z(_0192_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _8013_ (.A1(_1594_),
    .A2(_1622_),
    .ZN(_3132_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _8014_ (.A1(_0535_),
    .A2(_1295_),
    .B(_3132_),
    .ZN(_3133_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _8015_ (.A1(_0461_),
    .A2(_3120_),
    .ZN(_3134_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _8016_ (.A1(_3120_),
    .A2(_3133_),
    .B(_3134_),
    .ZN(_0193_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _8017_ (.A1(_0579_),
    .A2(_2399_),
    .ZN(_3135_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _8018_ (.I(_2794_),
    .Z(_3136_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _8019_ (.A1(_1558_),
    .A2(_3136_),
    .ZN(_3137_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _8020_ (.A1(_3135_),
    .A2(_3137_),
    .ZN(_3138_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _8021_ (.I0(_3138_),
    .I1(_0549_),
    .S(_3130_),
    .Z(_3139_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _8022_ (.I(_3139_),
    .Z(_0194_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _8023_ (.A1(_2736_),
    .A2(_3103_),
    .ZN(_3140_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _8024_ (.A1(_1290_),
    .A2(_3140_),
    .ZN(_3141_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _8025_ (.I0(_3141_),
    .I1(_0637_),
    .S(_3130_),
    .Z(_3142_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _8026_ (.I(_3142_),
    .Z(_0195_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _8027_ (.I(_1524_),
    .Z(_3143_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _8028_ (.I(_3143_),
    .Z(_3144_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _8029_ (.A1(_1706_),
    .A2(_1572_),
    .ZN(_3145_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _8030_ (.A1(_1530_),
    .A2(_3144_),
    .B(_3145_),
    .ZN(_3146_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _8031_ (.I0(_3146_),
    .I1(_0730_),
    .S(_3130_),
    .Z(_3147_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _8032_ (.I(_3147_),
    .Z(_0196_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _8033_ (.A1(_1710_),
    .A2(_1294_),
    .ZN(_3148_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _8034_ (.A1(_1626_),
    .A2(_3148_),
    .ZN(_3149_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _8035_ (.I0(_3149_),
    .I1(_0813_),
    .S(_3119_),
    .Z(_3150_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _8036_ (.I(_3150_),
    .Z(_0197_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _8037_ (.A1(_2416_),
    .A2(_1488_),
    .ZN(_0198_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _8038_ (.I(_3106_),
    .Z(_3151_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _8039_ (.A1(_3151_),
    .A2(_1677_),
    .ZN(_3152_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _8040_ (.I(_1685_),
    .Z(_3153_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _8041_ (.I(_2149_),
    .Z(_3154_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _8042_ (.A1(_2440_),
    .A2(_2461_),
    .ZN(_3155_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _8043_ (.A1(_1250_),
    .A2(_3155_),
    .ZN(_3156_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _8044_ (.I(_2503_),
    .Z(_3157_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _8045_ (.I(_3157_),
    .Z(_3158_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _8046_ (.A1(_1676_),
    .A2(_1268_),
    .ZN(_3159_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _8047_ (.A1(_3158_),
    .A2(_3159_),
    .ZN(_3160_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _8048_ (.A1(_3156_),
    .A2(_3160_),
    .B(_3059_),
    .ZN(_3161_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _8049_ (.A1(_1354_),
    .A2(_2348_),
    .ZN(_3162_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _8050_ (.I(_0898_),
    .Z(_3163_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _8051_ (.I(_3163_),
    .Z(_3164_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _8052_ (.A1(_2535_),
    .A2(_3162_),
    .B(_3164_),
    .ZN(_3165_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _8053_ (.A1(_1237_),
    .A2(_1045_),
    .A3(_1273_),
    .ZN(_3166_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_2 _8054_ (.A1(_1676_),
    .A2(_1236_),
    .A3(_1249_),
    .A4(_3166_),
    .ZN(_3167_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _8055_ (.A1(_3158_),
    .A2(_1370_),
    .B1(_3159_),
    .B2(_3167_),
    .ZN(_3168_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_2 _8056_ (.A1(_1612_),
    .A2(_1256_),
    .B(_1229_),
    .C(_2482_),
    .ZN(_3169_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _8057_ (.I(_3045_),
    .Z(_3170_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _8058_ (.A1(_1249_),
    .A2(_3159_),
    .B(_3169_),
    .C(_3170_),
    .ZN(_3171_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _8059_ (.A1(_3168_),
    .A2(_3171_),
    .ZN(_3172_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_1 _8060_ (.A1(_3154_),
    .A2(_3161_),
    .A3(_3165_),
    .B(_3172_),
    .ZN(_3173_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _8061_ (.A1(_1677_),
    .A2(_3153_),
    .B1(_2407_),
    .B2(_3173_),
    .ZN(_3174_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _8062_ (.I(_4241_),
    .Z(_3175_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _8063_ (.A1(_2618_),
    .A2(_0687_),
    .B(_2607_),
    .ZN(_3176_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _8064_ (.A1(_1354_),
    .A2(_3175_),
    .B(_2390_),
    .C(_3176_),
    .ZN(_3177_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _8065_ (.I(_1342_),
    .Z(_3178_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _8066_ (.A1(_0687_),
    .A2(_3175_),
    .ZN(_3179_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _8067_ (.A1(_3178_),
    .A2(_3179_),
    .ZN(_3180_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _8068_ (.I(_2384_),
    .Z(_3181_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _8069_ (.A1(_1272_),
    .A2(_3181_),
    .ZN(_3182_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _8070_ (.I(_3182_),
    .Z(_3183_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _8071_ (.I(_3183_),
    .Z(_3184_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _8072_ (.A1(_3177_),
    .A2(_3180_),
    .A3(_3184_),
    .ZN(_3185_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _8073_ (.A1(_4417_),
    .A2(_1279_),
    .ZN(_3186_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _8074_ (.A1(_2421_),
    .A2(_3186_),
    .ZN(_3187_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_1 _8075_ (.A1(_1570_),
    .A2(_3174_),
    .B1(_3185_),
    .B2(_3187_),
    .C(_2400_),
    .ZN(_3188_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _8076_ (.I(_1391_),
    .Z(_3189_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _8077_ (.A1(_3152_),
    .A2(_3188_),
    .B(_3189_),
    .ZN(_0199_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _8078_ (.A1(_3151_),
    .A2(_1678_),
    .ZN(_3190_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _8079_ (.I(_1498_),
    .Z(_3191_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _8080_ (.I(_2432_),
    .Z(_3192_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _8081_ (.A1(_3191_),
    .A2(_3192_),
    .B1(_3067_),
    .B2(_3154_),
    .ZN(_3193_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _8082_ (.I(_1685_),
    .Z(_3194_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _8083_ (.A1(_2383_),
    .A2(_3061_),
    .A3(_3192_),
    .ZN(_3195_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _8084_ (.A1(_3194_),
    .A2(_3156_),
    .B(_3195_),
    .ZN(_3196_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _8085_ (.A1(_3164_),
    .A2(_3196_),
    .ZN(_3197_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _8086_ (.A1(_2399_),
    .A2(_3167_),
    .ZN(_3198_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _8087_ (.I(_3170_),
    .Z(_3199_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _8088_ (.A1(_2383_),
    .A2(_3192_),
    .B(_3169_),
    .C(_3199_),
    .ZN(_3200_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _8089_ (.A1(_3193_),
    .A2(_3197_),
    .B1(_3198_),
    .B2(_3200_),
    .C(_2624_),
    .ZN(_3201_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _8090_ (.A1(_3178_),
    .A2(_3192_),
    .A3(_3179_),
    .ZN(_3202_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _8091_ (.A1(_2888_),
    .A2(_3202_),
    .ZN(_3203_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _8092_ (.A1(_3136_),
    .A2(_3061_),
    .A3(_3176_),
    .A4(_3203_),
    .ZN(_3204_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _8093_ (.A1(_3186_),
    .A2(_3204_),
    .B(_1576_),
    .ZN(_3205_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _8094_ (.A1(_3201_),
    .A2(_3205_),
    .B(_4201_),
    .ZN(_3206_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _8095_ (.A1(_3190_),
    .A2(_3206_),
    .B(_3189_),
    .ZN(_0200_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _8096_ (.I(_3106_),
    .Z(_3207_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _8097_ (.I(_3207_),
    .Z(_3208_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _8098_ (.I(_1348_),
    .Z(_3209_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _8099_ (.I(_3046_),
    .Z(_3210_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _8100_ (.A1(_2386_),
    .A2(_3090_),
    .B(_1370_),
    .ZN(_3211_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _8101_ (.A1(_3209_),
    .A2(_1507_),
    .Z(_3212_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _8102_ (.A1(_3090_),
    .A2(_1231_),
    .B(_3212_),
    .ZN(_3213_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _8103_ (.I(_3045_),
    .Z(_3214_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _8104_ (.A1(_1304_),
    .A2(_4175_),
    .B(_3214_),
    .ZN(_3215_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _8105_ (.I(_2388_),
    .Z(_3216_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _8106_ (.A1(_3211_),
    .A2(_3213_),
    .ZN(_3217_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_1 _8107_ (.A1(_3211_),
    .A2(_3213_),
    .B1(_3215_),
    .B2(_3216_),
    .C(_3217_),
    .ZN(_3218_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _8108_ (.I(_3158_),
    .Z(_3219_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _8109_ (.A1(_3219_),
    .A2(_3212_),
    .ZN(_3220_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _8110_ (.I(_2151_),
    .Z(_3221_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _8111_ (.A1(_3164_),
    .A2(_3221_),
    .B(_3067_),
    .ZN(_3222_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _8112_ (.A1(_4253_),
    .A2(_3153_),
    .B1(_2508_),
    .B2(_3059_),
    .C(_3191_),
    .ZN(_3223_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _8113_ (.A1(_3220_),
    .A2(_3222_),
    .B(_3223_),
    .ZN(_3224_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _8114_ (.A1(_3210_),
    .A2(_3218_),
    .A3(_3224_),
    .ZN(_3225_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _8115_ (.I(_1328_),
    .Z(_3226_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_1 _8116_ (.A1(_1429_),
    .A2(_1493_),
    .A3(_1494_),
    .B(_3220_),
    .ZN(_3227_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _8117_ (.A1(_3226_),
    .A2(_3227_),
    .B(_3207_),
    .ZN(_3228_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _8118_ (.I(_1301_),
    .Z(_3229_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _8119_ (.A1(_3208_),
    .A2(_3209_),
    .B1(_3225_),
    .B2(_3228_),
    .C(_3229_),
    .ZN(_0201_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _8120_ (.I(_3170_),
    .Z(_3230_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _8121_ (.A1(_1681_),
    .A2(_2155_),
    .B(_3221_),
    .ZN(_3231_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _8122_ (.A1(_3209_),
    .A2(_1507_),
    .ZN(_3232_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _8123_ (.A1(_0893_),
    .A2(_3232_),
    .Z(_3233_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _8124_ (.A1(_3230_),
    .A2(_3231_),
    .B(_3233_),
    .ZN(_3234_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _8125_ (.A1(_1451_),
    .A2(_3234_),
    .ZN(_3235_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _8126_ (.A1(_0869_),
    .A2(_2506_),
    .ZN(_3236_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _8127_ (.A1(_3081_),
    .A2(_3236_),
    .ZN(_3237_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _8128_ (.A1(_3179_),
    .A2(_3233_),
    .ZN(_3238_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _8129_ (.A1(_0687_),
    .A2(_2658_),
    .B1(_3178_),
    .B2(_3238_),
    .ZN(_3239_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _8130_ (.A1(_2624_),
    .A2(_3061_),
    .A3(_1339_),
    .A4(_2390_),
    .ZN(_3240_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _8131_ (.A1(_3239_),
    .A2(_3240_),
    .B(_4201_),
    .ZN(_3241_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _8132_ (.A1(_2633_),
    .A2(_3237_),
    .B(_3241_),
    .ZN(_3242_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _8133_ (.A1(_3151_),
    .A2(_0893_),
    .B1(_3235_),
    .B2(_3242_),
    .C(_3229_),
    .ZN(_0202_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _8134_ (.I(\as2650.cycle[4] ),
    .Z(_3243_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_4 _8135_ (.A1(_1486_),
    .A2(_0893_),
    .A3(_3209_),
    .A4(_1507_),
    .ZN(_3244_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _8136_ (.I(_1565_),
    .Z(_3245_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _8137_ (.A1(_3243_),
    .A2(_3244_),
    .B(_3245_),
    .ZN(_3246_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _8138_ (.A1(_3243_),
    .A2(_3244_),
    .B(_3246_),
    .ZN(_0203_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _8139_ (.A1(_3243_),
    .A2(_3244_),
    .ZN(_3247_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _8140_ (.A1(\as2650.cycle[5] ),
    .A2(_3247_),
    .Z(_3248_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _8141_ (.A1(_2416_),
    .A2(_3248_),
    .ZN(_0204_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _8142_ (.I(_1301_),
    .Z(_3249_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _8143_ (.I(_4171_),
    .Z(_3250_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _8144_ (.A1(_2150_),
    .A2(_3250_),
    .B(_1339_),
    .C(_3178_),
    .ZN(_3251_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_2 _8145_ (.A1(\as2650.cycle[5] ),
    .A2(_3243_),
    .A3(\as2650.cycle[3] ),
    .A4(_3232_),
    .ZN(_3252_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _8146_ (.A1(_2484_),
    .A2(_3252_),
    .Z(_3253_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _8147_ (.A1(_3175_),
    .A2(_3226_),
    .ZN(_3254_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _8148_ (.A1(_3226_),
    .A2(_3251_),
    .B1(_3253_),
    .B2(_3254_),
    .C(_3207_),
    .ZN(_3255_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _8149_ (.A1(_3208_),
    .A2(_2484_),
    .B(_3249_),
    .C(_3255_),
    .ZN(_0205_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _8150_ (.I(_2437_),
    .Z(_3256_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _8151_ (.I(_3256_),
    .Z(_3257_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_1 _8152_ (.A1(_1572_),
    .A2(_2477_),
    .A3(_2719_),
    .B(_3226_),
    .ZN(_3258_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _8153_ (.A1(_2484_),
    .A2(_3252_),
    .Z(_3259_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _8154_ (.A1(_1329_),
    .A2(_3259_),
    .Z(_3260_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _8155_ (.A1(_1570_),
    .A2(_3257_),
    .B1(_3258_),
    .B2(_3260_),
    .C(_3207_),
    .ZN(_3261_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _8156_ (.A1(_3208_),
    .A2(_1329_),
    .B(_3229_),
    .C(_3261_),
    .ZN(_0206_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _8157_ (.I(\as2650.psu[7] ),
    .ZN(_3262_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _8158_ (.I(net4),
    .ZN(_3263_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _8159_ (.A1(_3263_),
    .A2(_3074_),
    .A3(_1511_),
    .ZN(_3264_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _8160_ (.I(_4420_),
    .Z(_3265_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _8161_ (.A1(_3265_),
    .A2(_1527_),
    .ZN(_3266_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _8162_ (.A1(_1711_),
    .A2(_3266_),
    .ZN(_3267_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _8163_ (.A1(_4176_),
    .A2(_1510_),
    .ZN(_3268_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _8164_ (.A1(\as2650.psu[7] ),
    .A2(_2377_),
    .B(_3268_),
    .ZN(_3269_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _8165_ (.A1(_0791_),
    .A2(_3074_),
    .ZN(_3270_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _8166_ (.A1(_3267_),
    .A2(_3269_),
    .B(_3270_),
    .ZN(_3271_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _8167_ (.A1(_3264_),
    .A2(_3271_),
    .B(_3151_),
    .ZN(_3272_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _8168_ (.A1(_3262_),
    .A2(_3208_),
    .B(_3229_),
    .C(_3272_),
    .ZN(_0207_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_2 _8169_ (.A1(_0867_),
    .A2(_0879_),
    .A3(_1682_),
    .A4(_2346_),
    .ZN(_3273_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _8170_ (.A1(_3236_),
    .A2(_3273_),
    .ZN(_3274_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _8171_ (.A1(_2439_),
    .A2(_3186_),
    .ZN(_3275_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _8172_ (.A1(_0853_),
    .A2(_1248_),
    .A3(_2427_),
    .ZN(_3276_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _8173_ (.A1(_2428_),
    .A2(_3276_),
    .ZN(_3277_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _8174_ (.A1(_2631_),
    .A2(_3274_),
    .B(_3275_),
    .C(_3277_),
    .ZN(_3278_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _8175_ (.A1(_2336_),
    .A2(_0885_),
    .A3(_1462_),
    .ZN(_3279_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _8176_ (.A1(_2156_),
    .A2(_2506_),
    .B(_1364_),
    .C(_4200_),
    .ZN(_3280_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _8177_ (.A1(_1322_),
    .A2(_0889_),
    .B(_3279_),
    .C(_3280_),
    .ZN(_3281_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _8178_ (.A1(_1347_),
    .A2(_1363_),
    .Z(_3282_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_1 _8179_ (.A1(_4444_),
    .A2(_2435_),
    .A3(_3281_),
    .A4(_3282_),
    .ZN(_3283_));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _8180_ (.A1(_3073_),
    .A2(_3278_),
    .A3(_3283_),
    .Z(_3284_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_2 _8181_ (.A1(_3157_),
    .A2(_3163_),
    .A3(_1349_),
    .A4(_3065_),
    .ZN(_3285_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_2 _8182_ (.A1(_3052_),
    .A2(_3069_),
    .A3(_3071_),
    .ZN(_3286_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_2 _8183_ (.A1(_3055_),
    .A2(_3284_),
    .A3(_3285_),
    .A4(_3286_),
    .ZN(_3287_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _8184_ (.I(_3287_),
    .Z(_3288_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _8185_ (.I(_3288_),
    .Z(_3289_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _8186_ (.I(_1358_),
    .Z(_3290_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _8187_ (.I(_3290_),
    .Z(_3291_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _8188_ (.I(_3291_),
    .Z(_3292_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _8189_ (.I(_3095_),
    .Z(_3293_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _8190_ (.A1(_2144_),
    .A2(_1605_),
    .ZN(_3294_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _8191_ (.A1(_1544_),
    .A2(_2487_),
    .B(_3294_),
    .ZN(_3295_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _8192_ (.A1(_2144_),
    .A2(_1695_),
    .ZN(_3296_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _8193_ (.A1(_1695_),
    .A2(_3295_),
    .B(_3296_),
    .C(_1509_),
    .ZN(_3297_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _8194_ (.A1(_4392_),
    .A2(_2410_),
    .ZN(_3298_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _8195_ (.A1(_2899_),
    .A2(_2755_),
    .B(_1276_),
    .C(_3298_),
    .ZN(_3299_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _8196_ (.A1(_1442_),
    .A2(_3297_),
    .A3(_3299_),
    .ZN(_3300_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _8197_ (.A1(\as2650.pc[0] ),
    .A2(_4180_),
    .Z(_3301_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _8198_ (.A1(_3296_),
    .A2(_3301_),
    .Z(_3302_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_2 _8199_ (.A1(_2458_),
    .A2(_0834_),
    .A3(_2460_),
    .ZN(_3303_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _8200_ (.I0(_2145_),
    .I1(_3302_),
    .S(_3303_),
    .Z(_3304_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _8201_ (.A1(_2440_),
    .A2(_3302_),
    .ZN(_3305_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _8202_ (.A1(_0864_),
    .A2(_2440_),
    .B(_3305_),
    .C(_4161_),
    .ZN(_3306_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _8203_ (.A1(_4161_),
    .A2(_3304_),
    .B(_3306_),
    .C(_1251_),
    .ZN(_3307_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _8204_ (.A1(_3093_),
    .A2(_3300_),
    .A3(_3307_),
    .ZN(_3308_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _8205_ (.A1(_2754_),
    .A2(_4281_),
    .ZN(_3309_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _8206_ (.A1(_1549_),
    .A2(_3309_),
    .Z(_3310_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _8207_ (.A1(_2382_),
    .A2(_3310_),
    .ZN(_3311_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _8208_ (.A1(_0864_),
    .A2(_2854_),
    .B(_3058_),
    .C(_3311_),
    .ZN(_3312_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _8209_ (.A1(_3293_),
    .A2(_3308_),
    .A3(_3312_),
    .ZN(_3313_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _8210_ (.A1(_2335_),
    .A2(_3295_),
    .ZN(_3314_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _8211_ (.A1(_2145_),
    .A2(_2794_),
    .B(_3194_),
    .C(_3314_),
    .ZN(_3315_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _8212_ (.A1(_3214_),
    .A2(_3313_),
    .A3(_3315_),
    .ZN(_3316_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _8213_ (.I(_2387_),
    .Z(_3317_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _8214_ (.A1(\as2650.stack[7][0] ),
    .A2(_1919_),
    .B1(_1638_),
    .B2(\as2650.stack[6][0] ),
    .ZN(_3318_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _8215_ (.I(_1902_),
    .Z(_3319_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _8216_ (.I(_1654_),
    .Z(_3320_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_1 _8217_ (.A1(\as2650.stack[4][0] ),
    .A2(_3319_),
    .B1(_3320_),
    .B2(\as2650.stack[5][0] ),
    .C(_4475_),
    .ZN(_3321_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _8218_ (.I(_1637_),
    .Z(_3322_));
 gf180mcu_fd_sc_mcu7t5v0__oai222_1 _8219_ (.A1(\as2650.stack[3][0] ),
    .A2(_1918_),
    .B1(_1902_),
    .B2(\as2650.stack[0][0] ),
    .C1(\as2650.stack[1][0] ),
    .C2(_1654_),
    .ZN(_3323_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _8220_ (.I(_3323_),
    .ZN(_3324_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _8221_ (.A1(\as2650.stack[2][0] ),
    .A2(_3322_),
    .B(_0328_),
    .C(_3324_),
    .ZN(_3325_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _8222_ (.A1(_3318_),
    .A2(_3321_),
    .B(_3325_),
    .ZN(_3326_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _8223_ (.I(_2408_),
    .Z(_3327_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _8224_ (.A1(_0864_),
    .A2(_3317_),
    .B1(_3326_),
    .B2(_3327_),
    .ZN(_3328_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _8225_ (.I(_3290_),
    .Z(_3329_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _8226_ (.A1(_3316_),
    .A2(_3328_),
    .B(_3329_),
    .ZN(_3330_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _8227_ (.I(_3287_),
    .Z(_3331_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _8228_ (.A1(_0865_),
    .A2(_3292_),
    .B(_3330_),
    .C(_3331_),
    .ZN(_3332_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _8229_ (.A1(_0865_),
    .A2(_3289_),
    .B(_3332_),
    .C(_3112_),
    .ZN(_0208_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _8230_ (.I(_3291_),
    .Z(_3333_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _8231_ (.A1(_0910_),
    .A2(_2144_),
    .Z(_3334_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _8232_ (.I(_3334_),
    .Z(_3335_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _8233_ (.I(_2387_),
    .Z(_3336_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _8234_ (.A1(_3336_),
    .A2(_3335_),
    .ZN(_3337_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _8235_ (.A1(_1677_),
    .A2(_3335_),
    .B(_2926_),
    .ZN(_3338_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _8236_ (.A1(net6),
    .A2(_4281_),
    .ZN(_3339_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _8237_ (.A1(_4530_),
    .A2(_4380_),
    .A3(_3339_),
    .Z(_3340_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _8238_ (.A1(_4530_),
    .A2(_2503_),
    .ZN(_3341_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _8239_ (.A1(_2777_),
    .A2(_3340_),
    .B(_3341_),
    .C(_3089_),
    .ZN(_3342_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _8240_ (.A1(_1696_),
    .A2(_1681_),
    .A3(_3342_),
    .ZN(_3343_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _8241_ (.A1(_2362_),
    .A2(_3181_),
    .ZN(_3344_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _8242_ (.I(_2533_),
    .Z(_3345_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _8243_ (.A1(_4531_),
    .A2(_3345_),
    .ZN(_3346_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _8244_ (.A1(_3089_),
    .A2(_2438_),
    .A3(_3344_),
    .A4(_3346_),
    .ZN(_3347_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _8245_ (.A1(_1696_),
    .A2(_3334_),
    .B(_1276_),
    .ZN(_3348_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _8246_ (.A1(_1679_),
    .A2(_2545_),
    .ZN(_3349_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _8247_ (.A1(_0911_),
    .A2(_1618_),
    .B(_3349_),
    .ZN(_3350_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _8248_ (.A1(_3048_),
    .A2(_3348_),
    .B1(_3350_),
    .B2(_1696_),
    .ZN(_3351_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _8249_ (.A1(_2335_),
    .A2(_3347_),
    .A3(_3351_),
    .ZN(_3352_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _8250_ (.I(_3155_),
    .Z(_3353_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _8251_ (.A1(_1681_),
    .A2(_3353_),
    .ZN(_3354_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _8252_ (.A1(_0909_),
    .A2(_3301_),
    .Z(_3355_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _8253_ (.A1(_0911_),
    .A2(_3301_),
    .ZN(_3356_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _8254_ (.A1(_3355_),
    .A2(_3356_),
    .B(_3354_),
    .ZN(_3357_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _8255_ (.A1(_3354_),
    .A2(_3335_),
    .B(_3357_),
    .C(_1289_),
    .ZN(_3358_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _8256_ (.A1(_3338_),
    .A2(_3343_),
    .B(_3352_),
    .C(_3358_),
    .ZN(_3359_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _8257_ (.A1(\as2650.stack[3][1] ),
    .A2(_4474_),
    .B(_4473_),
    .ZN(_3360_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _8258_ (.I(_1903_),
    .Z(_3361_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _8259_ (.I(_1655_),
    .Z(_3362_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _8260_ (.A1(\as2650.stack[2][1] ),
    .A2(_1637_),
    .Z(_3363_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_1 _8261_ (.A1(\as2650.stack[0][1] ),
    .A2(_3361_),
    .B1(_3362_),
    .B2(\as2650.stack[1][1] ),
    .C(_3363_),
    .ZN(_3364_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _8262_ (.A1(\as2650.stack[4][1] ),
    .A2(_3361_),
    .B1(_3362_),
    .B2(\as2650.stack[5][1] ),
    .ZN(_3365_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _8263_ (.I(_1918_),
    .Z(_3366_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_1 _8264_ (.A1(\as2650.stack[7][1] ),
    .A2(_3366_),
    .B1(_3322_),
    .B2(\as2650.stack[6][1] ),
    .C(_4476_),
    .ZN(_3367_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _8265_ (.A1(_3360_),
    .A2(_3364_),
    .B1(_3365_),
    .B2(_3367_),
    .ZN(_3368_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _8266_ (.I(_2391_),
    .Z(_3369_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _8267_ (.A1(_3199_),
    .A2(_3359_),
    .B1(_3368_),
    .B2(_3369_),
    .ZN(_3370_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _8268_ (.I(_3290_),
    .Z(_3371_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _8269_ (.A1(_3337_),
    .A2(_3370_),
    .B(_3371_),
    .ZN(_3372_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _8270_ (.I(_3287_),
    .Z(_3373_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _8271_ (.I(_3373_),
    .Z(_3374_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _8272_ (.A1(_3333_),
    .A2(_3335_),
    .B(_3372_),
    .C(_3374_),
    .ZN(_3375_));
 gf180mcu_fd_sc_mcu7t5v0__and4_1 _8273_ (.A1(_3055_),
    .A2(_3284_),
    .A3(_3285_),
    .A4(_3286_),
    .Z(_3376_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _8274_ (.I(_3376_),
    .Z(_3377_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _8275_ (.A1(_2170_),
    .A2(_3377_),
    .B(_1566_),
    .ZN(_3378_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _8276_ (.A1(_3375_),
    .A2(_3378_),
    .ZN(_0209_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _8277_ (.I(_3291_),
    .Z(_3379_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _8278_ (.A1(_0910_),
    .A2(_0862_),
    .ZN(_3380_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _8279_ (.A1(_0919_),
    .A2(_3380_),
    .ZN(_3381_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _8280_ (.I(_3381_),
    .Z(_3382_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _8281_ (.A1(\as2650.stack[3][2] ),
    .A2(_4474_),
    .B(_4473_),
    .ZN(_3383_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _8282_ (.A1(\as2650.stack[2][2] ),
    .A2(_3322_),
    .ZN(_3384_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _8283_ (.A1(\as2650.stack[0][2] ),
    .A2(_3319_),
    .B1(_3320_),
    .B2(\as2650.stack[1][2] ),
    .ZN(_3385_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _8284_ (.I(_1637_),
    .Z(_3386_));
 gf180mcu_fd_sc_mcu7t5v0__oai222_1 _8285_ (.A1(\as2650.stack[7][2] ),
    .A2(_1918_),
    .B1(_1902_),
    .B2(\as2650.stack[4][2] ),
    .C1(\as2650.stack[5][2] ),
    .C2(_1654_),
    .ZN(_3387_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _8286_ (.A1(_0327_),
    .A2(_3387_),
    .ZN(_3388_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _8287_ (.A1(\as2650.stack[6][2] ),
    .A2(_3386_),
    .B(_3388_),
    .ZN(_3389_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_1 _8288_ (.A1(_3383_),
    .A2(_3384_),
    .A3(_3385_),
    .B(_3389_),
    .ZN(_3390_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _8289_ (.I(_3095_),
    .Z(_3391_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _8290_ (.A1(_1267_),
    .A2(_3057_),
    .B1(_3155_),
    .B2(_1288_),
    .ZN(_3392_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _8291_ (.I(_3392_),
    .Z(_3393_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_2 _8292_ (.A1(_1271_),
    .A2(_2157_),
    .A3(_3155_),
    .ZN(_3394_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _8293_ (.I(_3394_),
    .Z(_3395_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _8294_ (.A1(_0920_),
    .A2(_3355_),
    .ZN(_3396_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _8295_ (.A1(_3395_),
    .A2(_3396_),
    .ZN(_3397_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _8296_ (.A1(_3382_),
    .A2(_3393_),
    .B(_3397_),
    .ZN(_3398_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _8297_ (.A1(_0373_),
    .A2(_4517_),
    .ZN(_3399_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _8298_ (.A1(_1553_),
    .A2(_4517_),
    .Z(_3400_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _8299_ (.A1(_3399_),
    .A2(_3400_),
    .ZN(_3401_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _8300_ (.A1(_2581_),
    .A2(_4380_),
    .ZN(_3402_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _8301_ (.A1(_2581_),
    .A2(_4380_),
    .ZN(_3403_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _8302_ (.A1(_3339_),
    .A2(_3402_),
    .B(_3403_),
    .ZN(_3404_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _8303_ (.A1(_3401_),
    .A2(_3404_),
    .Z(_3405_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _8304_ (.A1(_1553_),
    .A2(_2538_),
    .ZN(_3406_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _8305_ (.A1(_2509_),
    .A2(_3405_),
    .B(_3406_),
    .ZN(_3407_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _8306_ (.A1(_0919_),
    .A2(_1708_),
    .ZN(_3408_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _8307_ (.A1(_1336_),
    .A2(_2620_),
    .B(_3408_),
    .ZN(_3409_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _8308_ (.A1(_2365_),
    .A2(_2754_),
    .ZN(_3410_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _8309_ (.A1(_0376_),
    .A2(_2533_),
    .B(_1508_),
    .C(_3410_),
    .ZN(_3411_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _8310_ (.A1(_3082_),
    .A2(_3381_),
    .B1(_3409_),
    .B2(_2645_),
    .C(_3411_),
    .ZN(_3412_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _8311_ (.A1(_3093_),
    .A2(_3412_),
    .ZN(_3413_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _8312_ (.A1(_3070_),
    .A2(_3407_),
    .B(_3413_),
    .ZN(_3414_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _8313_ (.I(_2437_),
    .Z(_3415_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _8314_ (.A1(_3415_),
    .A2(_3382_),
    .B1(_3409_),
    .B2(_2549_),
    .C(_2856_),
    .ZN(_3416_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _8315_ (.A1(_3391_),
    .A2(_3398_),
    .B1(_3414_),
    .B2(_2345_),
    .C(_3416_),
    .ZN(_3417_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _8316_ (.A1(_3336_),
    .A2(_3382_),
    .B1(_3390_),
    .B2(_3369_),
    .C(_3417_),
    .ZN(_3418_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _8317_ (.A1(_3329_),
    .A2(_3382_),
    .ZN(_3419_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _8318_ (.I(_3376_),
    .Z(_3420_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _8319_ (.A1(_3379_),
    .A2(_3418_),
    .B(_3419_),
    .C(_3420_),
    .ZN(_3421_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _8320_ (.A1(_2178_),
    .A2(_3377_),
    .B(_3421_),
    .ZN(_3422_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _8321_ (.A1(_2416_),
    .A2(_3422_),
    .ZN(_0210_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _8322_ (.A1(\as2650.pc[2] ),
    .A2(_0909_),
    .A3(\as2650.pc[0] ),
    .ZN(_3423_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _8323_ (.A1(_0927_),
    .A2(_3423_),
    .Z(_3424_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _8324_ (.I(_3424_),
    .Z(_3425_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _8325_ (.I(_2387_),
    .Z(_3426_));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _8326_ (.A1(_2181_),
    .A2(_0919_),
    .A3(_3355_),
    .Z(_3427_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _8327_ (.I(_3427_),
    .Z(_3428_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _8328_ (.A1(_0920_),
    .A2(_3355_),
    .B(_2182_),
    .ZN(_3429_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _8329_ (.A1(_1293_),
    .A2(_3353_),
    .ZN(_3430_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _8330_ (.A1(_3428_),
    .A2(_3429_),
    .B(_3430_),
    .ZN(_3431_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _8331_ (.A1(_2182_),
    .A2(_1617_),
    .ZN(_3432_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _8332_ (.A1(_1708_),
    .A2(_2641_),
    .B(_3432_),
    .ZN(_3433_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _8333_ (.A1(_2368_),
    .A2(_1490_),
    .B(_1508_),
    .C(_2651_),
    .ZN(_3434_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _8334_ (.A1(_2494_),
    .A2(_3424_),
    .B1(_3433_),
    .B2(_2352_),
    .C(_3434_),
    .ZN(_3435_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _8335_ (.A1(_2793_),
    .A2(_3435_),
    .B(_3076_),
    .ZN(_3436_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _8336_ (.A1(_3156_),
    .A2(_3425_),
    .B(_3431_),
    .C(_3436_),
    .ZN(_3437_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _8337_ (.I(_3399_),
    .ZN(_3438_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _8338_ (.A1(_3400_),
    .A2(_3404_),
    .B(_3438_),
    .ZN(_3439_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _8339_ (.A1(_0508_),
    .A2(_0366_),
    .A3(_3439_),
    .Z(_3440_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _8340_ (.A1(_1147_),
    .A2(_3157_),
    .ZN(_3441_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _8341_ (.A1(_3181_),
    .A2(_3440_),
    .B(_3441_),
    .C(_2925_),
    .ZN(_3442_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _8342_ (.A1(_2854_),
    .A2(_3425_),
    .B(_3442_),
    .C(_3058_),
    .ZN(_3443_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _8343_ (.A1(_3293_),
    .A2(_3437_),
    .A3(_3443_),
    .ZN(_3444_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _8344_ (.A1(_3415_),
    .A2(_3424_),
    .B1(_3433_),
    .B2(_2524_),
    .C(_2856_),
    .ZN(_3445_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _8345_ (.I(_3445_),
    .ZN(_3446_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _8346_ (.A1(\as2650.stack[3][3] ),
    .A2(_1919_),
    .B1(_1638_),
    .B2(\as2650.stack[2][3] ),
    .ZN(_3447_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_1 _8347_ (.A1(\as2650.stack[0][3] ),
    .A2(_1903_),
    .B1(_1655_),
    .B2(\as2650.stack[1][3] ),
    .C(_0328_),
    .ZN(_3448_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _8348_ (.A1(\as2650.stack[4][3] ),
    .A2(_1903_),
    .B1(_1655_),
    .B2(\as2650.stack[5][3] ),
    .ZN(_3449_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_1 _8349_ (.A1(\as2650.stack[7][3] ),
    .A2(_1919_),
    .B1(_1638_),
    .B2(\as2650.stack[6][3] ),
    .C(_4475_),
    .ZN(_3450_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _8350_ (.A1(_3447_),
    .A2(_3448_),
    .B1(_3449_),
    .B2(_3450_),
    .ZN(_3451_));
 gf180mcu_fd_sc_mcu7t5v0__aoi222_1 _8351_ (.A1(_3426_),
    .A2(_3425_),
    .B1(_3444_),
    .B2(_3446_),
    .C1(_3451_),
    .C2(_3327_),
    .ZN(_3452_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _8352_ (.A1(_3371_),
    .A2(_3452_),
    .B(_3420_),
    .ZN(_3453_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _8353_ (.A1(_3333_),
    .A2(_3425_),
    .B(_3453_),
    .ZN(_3454_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _8354_ (.A1(_0928_),
    .A2(_3289_),
    .B(_3454_),
    .C(_3112_),
    .ZN(_0211_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _8355_ (.A1(_0927_),
    .A2(_3423_),
    .ZN(_3455_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _8356_ (.A1(_2188_),
    .A2(_3455_),
    .Z(_3456_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _8357_ (.I(_3456_),
    .Z(_3457_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _8358_ (.I(_3393_),
    .Z(_3458_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _8359_ (.I(_3394_),
    .Z(_3459_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _8360_ (.A1(_2189_),
    .A2(_3428_),
    .ZN(_3460_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _8361_ (.A1(_2189_),
    .A2(_3428_),
    .Z(_3461_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _8362_ (.A1(_3460_),
    .A2(_3461_),
    .B(_1685_),
    .ZN(_3462_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _8363_ (.A1(_2188_),
    .A2(_1605_),
    .ZN(_3463_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _8364_ (.A1(_1679_),
    .A2(_2698_),
    .B(_3463_),
    .ZN(_3464_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _8365_ (.A1(_3256_),
    .A2(_3457_),
    .B1(_3464_),
    .B2(_2524_),
    .C(_2927_),
    .ZN(_3465_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _8366_ (.A1(_0506_),
    .A2(_0366_),
    .ZN(_3466_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _8367_ (.A1(_0506_),
    .A2(_0366_),
    .ZN(_3467_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _8368_ (.A1(_3466_),
    .A2(_3439_),
    .B(_3467_),
    .ZN(_3468_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _8369_ (.A1(_1581_),
    .A2(_0496_),
    .A3(_3468_),
    .Z(_3469_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _8370_ (.A1(_0596_),
    .A2(_1490_),
    .ZN(_3470_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _8371_ (.A1(_1267_),
    .A2(_0898_),
    .ZN(_3471_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _8372_ (.A1(_2648_),
    .A2(_3469_),
    .B(_3470_),
    .C(_3471_),
    .ZN(_3472_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _8373_ (.A1(_2353_),
    .A2(_3464_),
    .ZN(_3473_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _8374_ (.A1(\as2650.addr_buff[4] ),
    .A2(_2754_),
    .ZN(_3474_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_2 _8375_ (.A1(_1582_),
    .A2(_2533_),
    .B(_1508_),
    .C(_3474_),
    .ZN(_3475_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _8376_ (.A1(_3082_),
    .A2(_3456_),
    .B(_3475_),
    .ZN(_3476_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _8377_ (.A1(_2482_),
    .A2(_2354_),
    .A3(_3473_),
    .A4(_3476_),
    .ZN(_3477_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _8378_ (.A1(_3472_),
    .A2(_3477_),
    .ZN(_3478_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _8379_ (.A1(_3459_),
    .A2(_3462_),
    .B(_3465_),
    .C(_3478_),
    .ZN(_3479_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _8380_ (.A1(_3458_),
    .A2(_3457_),
    .B1(_3479_),
    .B2(_3291_),
    .ZN(_3480_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _8381_ (.I(_2391_),
    .Z(_3481_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _8382_ (.A1(\as2650.stack[3][4] ),
    .A2(_2215_),
    .B(_4473_),
    .ZN(_3482_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _8383_ (.A1(\as2650.stack[2][4] ),
    .A2(_1639_),
    .ZN(_3483_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _8384_ (.A1(\as2650.stack[0][4] ),
    .A2(_1904_),
    .B1(_1656_),
    .B2(\as2650.stack[1][4] ),
    .ZN(_3484_));
 gf180mcu_fd_sc_mcu7t5v0__oai222_1 _8385_ (.A1(\as2650.stack[4][4] ),
    .A2(_3319_),
    .B1(_3322_),
    .B2(\as2650.stack[6][4] ),
    .C1(_3320_),
    .C2(\as2650.stack[5][4] ),
    .ZN(_3485_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _8386_ (.A1(_0525_),
    .A2(_3485_),
    .ZN(_3486_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _8387_ (.A1(\as2650.stack[7][4] ),
    .A2(_1920_),
    .B(_3486_),
    .ZN(_3487_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_1 _8388_ (.A1(_3482_),
    .A2(_3483_),
    .A3(_3484_),
    .B(_3487_),
    .ZN(_3488_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _8389_ (.A1(_3481_),
    .A2(_3488_),
    .ZN(_3489_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _8390_ (.A1(_3480_),
    .A2(_3489_),
    .ZN(_3490_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _8391_ (.A1(_3210_),
    .A2(_3457_),
    .B(_3490_),
    .ZN(_3491_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _8392_ (.I(_2388_),
    .Z(_3492_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _8393_ (.A1(_3492_),
    .A2(_3457_),
    .B(_3288_),
    .ZN(_3493_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _8394_ (.A1(_0933_),
    .A2(_3374_),
    .B1(_3491_),
    .B2(_3493_),
    .C(_2415_),
    .ZN(_0212_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_2 _8395_ (.A1(_0933_),
    .A2(_0927_),
    .A3(_3423_),
    .ZN(_3494_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _8396_ (.A1(_2195_),
    .A2(_3494_),
    .Z(_3495_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _8397_ (.I(_3495_),
    .ZN(_3496_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _8398_ (.A1(_3393_),
    .A2(_3496_),
    .ZN(_3497_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _8399_ (.A1(_1579_),
    .A2(_2762_),
    .ZN(_3498_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _8400_ (.A1(_0939_),
    .A2(_1614_),
    .B(_3498_),
    .ZN(_3499_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _8401_ (.A1(_4265_),
    .A2(_3157_),
    .ZN(_3500_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _8402_ (.A1(_0685_),
    .A2(_2539_),
    .B(_2396_),
    .ZN(_3501_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _8403_ (.A1(_2996_),
    .A2(_3496_),
    .B1(_3500_),
    .B2(_3501_),
    .ZN(_3502_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _8404_ (.A1(_3221_),
    .A2(_3499_),
    .B(_3502_),
    .C(_1294_),
    .ZN(_3503_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _8405_ (.I(_3471_),
    .Z(_3504_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _8406_ (.A1(_2694_),
    .A2(_0496_),
    .Z(_3505_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _8407_ (.A1(_2694_),
    .A2(_0496_),
    .Z(_3506_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _8408_ (.A1(_3505_),
    .A2(_3468_),
    .B(_3506_),
    .ZN(_3507_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _8409_ (.A1(_1180_),
    .A2(_0583_),
    .A3(_3507_),
    .Z(_3508_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _8410_ (.A1(_2509_),
    .A2(_3508_),
    .ZN(_3509_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _8411_ (.A1(_2736_),
    .A2(_2756_),
    .B(_3504_),
    .C(_3509_),
    .ZN(_3510_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _8412_ (.A1(_2196_),
    .A2(_2189_),
    .A3(_3428_),
    .ZN(_3511_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _8413_ (.A1(_0940_),
    .A2(_3460_),
    .ZN(_3512_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _8414_ (.A1(_3395_),
    .A2(_3511_),
    .A3(_3512_),
    .ZN(_3513_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _8415_ (.A1(_3059_),
    .A2(_3503_),
    .B(_3510_),
    .C(_3513_),
    .ZN(_3514_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _8416_ (.A1(_3497_),
    .A2(_3514_),
    .B(_3391_),
    .ZN(_3515_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_1 _8417_ (.A1(_3250_),
    .A2(_3495_),
    .B1(_3499_),
    .B2(_2513_),
    .C(_3154_),
    .ZN(_3516_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _8418_ (.A1(_3515_),
    .A2(_3516_),
    .ZN(_3517_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _8419_ (.I(\as2650.stack[2][5] ),
    .ZN(_3518_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _8420_ (.A1(\as2650.stack[3][5] ),
    .A2(_2215_),
    .ZN(_3519_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _8421_ (.A1(\as2650.stack[0][5] ),
    .A2(_3361_),
    .B1(_3362_),
    .B2(\as2650.stack[1][5] ),
    .ZN(_3520_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _8422_ (.A1(_3518_),
    .A2(_0426_),
    .B1(_3519_),
    .B2(_4453_),
    .C(_3520_),
    .ZN(_3521_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _8423_ (.A1(\as2650.stack[7][5] ),
    .A2(_3366_),
    .B1(_3386_),
    .B2(\as2650.stack[6][5] ),
    .ZN(_3522_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _8424_ (.A1(\as2650.stack[4][5] ),
    .A2(_1904_),
    .B1(_1656_),
    .B2(\as2650.stack[5][5] ),
    .ZN(_3523_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _8425_ (.A1(_0525_),
    .A2(_3522_),
    .A3(_3523_),
    .ZN(_3524_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _8426_ (.A1(_3521_),
    .A2(_3524_),
    .ZN(_3525_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _8427_ (.I(_3290_),
    .Z(_3526_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _8428_ (.A1(_3336_),
    .A2(_3496_),
    .B1(_3525_),
    .B2(_3369_),
    .C(_3526_),
    .ZN(_3527_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _8429_ (.A1(_3379_),
    .A2(_3495_),
    .B1(_3517_),
    .B2(_3527_),
    .C(_3373_),
    .ZN(_3528_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _8430_ (.A1(_0940_),
    .A2(_3289_),
    .B(_3528_),
    .C(_3112_),
    .ZN(_0213_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _8431_ (.A1(_2195_),
    .A2(_3494_),
    .ZN(_3529_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _8432_ (.A1(_0946_),
    .A2(_3529_),
    .ZN(_3530_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _8433_ (.A1(_0946_),
    .A2(_1618_),
    .ZN(_3531_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _8434_ (.A1(_1709_),
    .A2(_2790_),
    .B(_3531_),
    .ZN(_3532_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _8435_ (.I(_2645_),
    .Z(_3533_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _8436_ (.A1(_0759_),
    .A2(_2539_),
    .ZN(_3534_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _8437_ (.A1(_4357_),
    .A2(_3345_),
    .B(_3534_),
    .ZN(_3535_));
 gf180mcu_fd_sc_mcu7t5v0__aoi222_1 _8438_ (.A1(_2495_),
    .A2(_3530_),
    .B1(_3532_),
    .B2(_3533_),
    .C1(_3089_),
    .C2(_3535_),
    .ZN(_3536_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _8439_ (.A1(_0758_),
    .A2(_0674_),
    .Z(_3537_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _8440_ (.A1(_2800_),
    .A2(_0583_),
    .ZN(_3538_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _8441_ (.A1(_2800_),
    .A2(_0583_),
    .ZN(_3539_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _8442_ (.A1(_3538_),
    .A2(_3507_),
    .B(_3539_),
    .ZN(_3540_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _8443_ (.A1(_3537_),
    .A2(_3540_),
    .Z(_3541_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _8444_ (.A1(_3537_),
    .A2(_3540_),
    .B(_3181_),
    .ZN(_3542_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_2 _8445_ (.A1(_1526_),
    .A2(_2777_),
    .B1(_3541_),
    .B2(_3542_),
    .C(_3070_),
    .ZN(_3543_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _8446_ (.A1(_3164_),
    .A2(_3536_),
    .B(_3543_),
    .ZN(_3544_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _8447_ (.A1(_0946_),
    .A2(_3511_),
    .Z(_3545_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _8448_ (.A1(_3459_),
    .A2(_3545_),
    .ZN(_3546_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_1 _8449_ (.A1(_3458_),
    .A2(_3530_),
    .B1(_3544_),
    .B2(_3126_),
    .C(_3546_),
    .ZN(_3547_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_1 _8450_ (.A1(_3250_),
    .A2(_3530_),
    .B1(_3532_),
    .B2(_2513_),
    .C(_3154_),
    .ZN(_3548_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _8451_ (.A1(_3153_),
    .A2(_3547_),
    .B(_3548_),
    .ZN(_3549_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _8452_ (.A1(_0947_),
    .A2(_3529_),
    .Z(_3550_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _8453_ (.A1(\as2650.stack[0][6] ),
    .A2(_3319_),
    .B1(_3320_),
    .B2(\as2650.stack[1][6] ),
    .ZN(_3551_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _8454_ (.I(_3551_),
    .ZN(_3552_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_1 _8455_ (.A1(\as2650.stack[3][6] ),
    .A2(_1920_),
    .B1(_3386_),
    .B2(\as2650.stack[2][6] ),
    .C(_3552_),
    .ZN(_3553_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _8456_ (.A1(\as2650.stack[7][6] ),
    .A2(_3366_),
    .B1(_3386_),
    .B2(\as2650.stack[6][6] ),
    .ZN(_3554_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_1 _8457_ (.A1(\as2650.stack[4][6] ),
    .A2(_1904_),
    .B1(_1656_),
    .B2(\as2650.stack[5][6] ),
    .C(_4476_),
    .ZN(_3555_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _8458_ (.A1(_4477_),
    .A2(_3553_),
    .B1(_3554_),
    .B2(_3555_),
    .ZN(_3556_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _8459_ (.I(_3556_),
    .ZN(_3557_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _8460_ (.A1(_3216_),
    .A2(_3550_),
    .B1(_3557_),
    .B2(_3481_),
    .C(_3371_),
    .ZN(_3558_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _8461_ (.A1(_3333_),
    .A2(_3530_),
    .B1(_3549_),
    .B2(_3558_),
    .C(_3288_),
    .ZN(_3559_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _8462_ (.A1(_2201_),
    .A2(_3377_),
    .B(_1566_),
    .ZN(_3560_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _8463_ (.A1(_3559_),
    .A2(_3560_),
    .ZN(_0214_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _8464_ (.A1(_0945_),
    .A2(_2194_),
    .A3(_3494_),
    .ZN(_3561_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _8465_ (.A1(_0953_),
    .A2(_3561_),
    .Z(_3562_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _8466_ (.I(_3562_),
    .Z(_3563_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _8467_ (.A1(_2825_),
    .A2(_0674_),
    .Z(_3564_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _8468_ (.A1(_2825_),
    .A2(_0674_),
    .Z(_3565_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _8469_ (.A1(_3564_),
    .A2(_3540_),
    .B(_3565_),
    .ZN(_3566_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _8470_ (.A1(_1604_),
    .A2(_4370_),
    .A3(_3566_),
    .Z(_3567_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _8471_ (.A1(_3345_),
    .A2(_3567_),
    .ZN(_3568_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _8472_ (.A1(_1619_),
    .A2(_2540_),
    .B(_3504_),
    .C(_3568_),
    .ZN(_3569_));
 gf180mcu_fd_sc_mcu7t5v0__and4_1 _8473_ (.A1(_0945_),
    .A2(_2195_),
    .A3(_2187_),
    .A4(_3427_),
    .Z(_3570_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _8474_ (.A1(_2203_),
    .A2(_3570_),
    .Z(_3571_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _8475_ (.A1(_2925_),
    .A2(_3163_),
    .B(_3156_),
    .ZN(_3572_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _8476_ (.A1(_0953_),
    .A2(_1605_),
    .ZN(_3573_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _8477_ (.A1(_1679_),
    .A2(_2849_),
    .B(_3573_),
    .ZN(_3574_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _8478_ (.A1(_2153_),
    .A2(_1489_),
    .ZN(_3575_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _8479_ (.A1(_1599_),
    .A2(_1490_),
    .B(_3575_),
    .ZN(_3576_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_1 _8480_ (.A1(_2526_),
    .A2(_3562_),
    .B1(_3576_),
    .B2(_1509_),
    .C(_2481_),
    .ZN(_3577_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _8481_ (.A1(_2645_),
    .A2(_3574_),
    .B(_3577_),
    .C(_3076_),
    .ZN(_3578_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _8482_ (.A1(_3395_),
    .A2(_3571_),
    .B1(_3563_),
    .B2(_3572_),
    .C(_3578_),
    .ZN(_3579_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _8483_ (.A1(_3293_),
    .A2(_3569_),
    .A3(_3579_),
    .ZN(_3580_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _8484_ (.A1(_3415_),
    .A2(_3563_),
    .ZN(_3581_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _8485_ (.A1(_2492_),
    .A2(_3574_),
    .B(_3581_),
    .C(_3001_),
    .ZN(_3582_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _8486_ (.A1(\as2650.stack[3][7] ),
    .A2(_1920_),
    .B1(_1639_),
    .B2(\as2650.stack[2][7] ),
    .ZN(_3583_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_1 _8487_ (.A1(\as2650.stack[0][7] ),
    .A2(_1905_),
    .B1(_1657_),
    .B2(\as2650.stack[1][7] ),
    .C(_0525_),
    .ZN(_3584_));
 gf180mcu_fd_sc_mcu7t5v0__oai222_1 _8488_ (.A1(\as2650.stack[7][7] ),
    .A2(_3366_),
    .B1(_3361_),
    .B2(\as2650.stack[4][7] ),
    .C1(\as2650.stack[5][7] ),
    .C2(_3362_),
    .ZN(_3585_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _8489_ (.I(_3585_),
    .ZN(_3586_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _8490_ (.A1(\as2650.stack[6][7] ),
    .A2(_1639_),
    .B(_4476_),
    .C(_3586_),
    .ZN(_3587_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _8491_ (.A1(_3583_),
    .A2(_3584_),
    .B(_3587_),
    .ZN(_3588_));
 gf180mcu_fd_sc_mcu7t5v0__aoi222_1 _8492_ (.A1(_3317_),
    .A2(_3563_),
    .B1(_3580_),
    .B2(_3582_),
    .C1(_3588_),
    .C2(_2391_),
    .ZN(_3589_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _8493_ (.A1(_3371_),
    .A2(_3589_),
    .B(_3376_),
    .ZN(_3590_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _8494_ (.A1(_3333_),
    .A2(_3563_),
    .B(_3590_),
    .ZN(_3591_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _8495_ (.I(_2577_),
    .Z(_3592_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _8496_ (.A1(_0953_),
    .A2(_3289_),
    .B(_3591_),
    .C(_3592_),
    .ZN(_0215_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _8497_ (.A1(_0966_),
    .A2(_3374_),
    .ZN(_3593_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _8498_ (.A1(_0952_),
    .A2(_3561_),
    .ZN(_3594_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _8499_ (.A1(_0965_),
    .A2(_3594_),
    .Z(_3595_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _8500_ (.I(_3595_),
    .Z(_3596_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _8501_ (.A1(\as2650.pc[8] ),
    .A2(_2203_),
    .A3(_3570_),
    .ZN(_3597_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _8502_ (.I(_3057_),
    .Z(_3598_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _8503_ (.A1(_2204_),
    .A2(_3570_),
    .B(_0965_),
    .ZN(_3599_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_1 _8504_ (.A1(_3103_),
    .A2(_3598_),
    .A3(_3353_),
    .A4(_3599_),
    .ZN(_3600_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _8505_ (.A1(_0965_),
    .A2(_1618_),
    .ZN(_3601_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _8506_ (.A1(_1709_),
    .A2(_2903_),
    .B(_3601_),
    .ZN(_3602_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _8507_ (.A1(_1549_),
    .A2(_2539_),
    .ZN(_3603_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _8508_ (.A1(_2334_),
    .A2(_2755_),
    .B(_1509_),
    .C(_3603_),
    .ZN(_3604_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _8509_ (.A1(_2996_),
    .A2(_3595_),
    .Z(_3605_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _8510_ (.A1(_3533_),
    .A2(_3602_),
    .B(_3604_),
    .C(_3605_),
    .ZN(_3606_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _8511_ (.A1(_1616_),
    .A2(_4370_),
    .ZN(_3607_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _8512_ (.A1(_1616_),
    .A2(_4370_),
    .ZN(_3608_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _8513_ (.A1(_3607_),
    .A2(_3566_),
    .B(_3608_),
    .ZN(_3609_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _8514_ (.A1(_0896_),
    .A2(_3609_),
    .ZN(_3610_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _8515_ (.A1(_2899_),
    .A2(_3610_),
    .Z(_3611_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _8516_ (.A1(_3598_),
    .A2(_3606_),
    .B1(_3611_),
    .B2(_3070_),
    .ZN(_3612_));
 gf180mcu_fd_sc_mcu7t5v0__aoi222_1 _8517_ (.A1(_3597_),
    .A2(_3600_),
    .B1(_3596_),
    .B2(_3572_),
    .C1(_1443_),
    .C2(_3612_),
    .ZN(_3613_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _8518_ (.A1(_3257_),
    .A2(_3596_),
    .B1(_3602_),
    .B2(_2550_),
    .C(_2928_),
    .ZN(_3614_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _8519_ (.A1(_3391_),
    .A2(_3613_),
    .B(_3614_),
    .ZN(_3615_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _8520_ (.A1(_3426_),
    .A2(_3596_),
    .ZN(_3616_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _8521_ (.A1(_1085_),
    .A2(_1499_),
    .B(_3046_),
    .C(_3616_),
    .ZN(_3617_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_1 _8522_ (.A1(_3210_),
    .A2(_3596_),
    .B1(_3615_),
    .B2(_3617_),
    .C(_3420_),
    .ZN(_3618_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _8523_ (.I(_1391_),
    .Z(_3619_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _8524_ (.A1(_3593_),
    .A2(_3618_),
    .B(_3619_),
    .ZN(_0216_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _8525_ (.I(_2911_),
    .Z(_3620_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _8526_ (.I(_3288_),
    .Z(_3621_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _8527_ (.A1(_0964_),
    .A2(_3594_),
    .ZN(_3622_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _8528_ (.A1(_3620_),
    .A2(_3622_),
    .Z(_3623_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _8529_ (.I(_3623_),
    .Z(_3624_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _8530_ (.A1(_2382_),
    .A2(_3058_),
    .ZN(_3625_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _8531_ (.A1(_2333_),
    .A2(_3610_),
    .ZN(_3626_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _8532_ (.A1(_2362_),
    .A2(_3626_),
    .ZN(_3627_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _8533_ (.A1(_3620_),
    .A2(_3597_),
    .Z(_3628_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _8534_ (.A1(_0979_),
    .A2(_1708_),
    .ZN(_3629_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _8535_ (.A1(_1336_),
    .A2(_2936_),
    .B(_3629_),
    .ZN(_3630_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _8536_ (.A1(_3221_),
    .A2(_3630_),
    .ZN(_3631_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _8537_ (.A1(\as2650.addr_buff[1] ),
    .A2(_2538_),
    .ZN(_3632_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _8538_ (.A1(_1275_),
    .A2(_3341_),
    .A3(_3632_),
    .ZN(_3633_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _8539_ (.A1(_2526_),
    .A2(_3623_),
    .B(_3633_),
    .C(_1234_),
    .ZN(_3634_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_1 _8540_ (.A1(_3076_),
    .A2(_3631_),
    .A3(_3634_),
    .B(_3095_),
    .ZN(_3635_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _8541_ (.A1(_3572_),
    .A2(_3624_),
    .B1(_3628_),
    .B2(_3395_),
    .C(_3635_),
    .ZN(_3636_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _8542_ (.A1(_3625_),
    .A2(_3627_),
    .B(_3636_),
    .ZN(_3637_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _8543_ (.A1(_3257_),
    .A2(_3624_),
    .B1(_3630_),
    .B2(_2549_),
    .C(_2928_),
    .ZN(_3638_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _8544_ (.I(_3638_),
    .ZN(_3639_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _8545_ (.A1(_3637_),
    .A2(_3639_),
    .ZN(_3640_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _8546_ (.A1(_0335_),
    .A2(_3369_),
    .B1(_3317_),
    .B2(_3624_),
    .ZN(_3641_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _8547_ (.A1(_3640_),
    .A2(_3641_),
    .B(_3329_),
    .ZN(_3642_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _8548_ (.A1(_3292_),
    .A2(_3624_),
    .B(_3642_),
    .C(_3331_),
    .ZN(_3643_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _8549_ (.A1(_3620_),
    .A2(_3621_),
    .B(_3643_),
    .C(_3592_),
    .ZN(_0217_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _8550_ (.A1(\as2650.pc[9] ),
    .A2(\as2650.pc[8] ),
    .A3(_3594_),
    .ZN(_3644_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _8551_ (.A1(_2969_),
    .A2(_3644_),
    .Z(_3645_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _8552_ (.A1(_2952_),
    .A2(_3610_),
    .ZN(_3646_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _8553_ (.A1(_2365_),
    .A2(_3646_),
    .ZN(_3647_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _8554_ (.A1(_3620_),
    .A2(_3597_),
    .ZN(_3648_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _8555_ (.A1(_2969_),
    .A2(_3648_),
    .Z(_3649_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _8556_ (.A1(_0990_),
    .A2(_1544_),
    .ZN(_3650_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _8557_ (.A1(_1709_),
    .A2(_2976_),
    .B(_3650_),
    .ZN(_3651_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _8558_ (.A1(_0989_),
    .A2(_3644_),
    .Z(_3652_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _8559_ (.A1(_2395_),
    .A2(_3406_),
    .ZN(_3653_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _8560_ (.A1(_2365_),
    .A2(_2776_),
    .B(_3653_),
    .ZN(_3654_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _8561_ (.A1(_2527_),
    .A2(_3652_),
    .B(_3654_),
    .C(_2160_),
    .ZN(_3655_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _8562_ (.A1(_3533_),
    .A2(_3651_),
    .B(_3655_),
    .ZN(_3656_));
 gf180mcu_fd_sc_mcu7t5v0__aoi222_1 _8563_ (.A1(_3504_),
    .A2(_3647_),
    .B1(_3649_),
    .B2(_3459_),
    .C1(_3103_),
    .C2(_3656_),
    .ZN(_3657_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _8564_ (.A1(_3458_),
    .A2(_3645_),
    .B(_3657_),
    .C(_3391_),
    .ZN(_3658_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_1 _8565_ (.A1(_3250_),
    .A2(_3645_),
    .B1(_3651_),
    .B2(_2492_),
    .C(_3001_),
    .ZN(_3659_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _8566_ (.A1(_3658_),
    .A2(_3659_),
    .ZN(_3660_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _8567_ (.A1(_0436_),
    .A2(_3481_),
    .B1(_3426_),
    .B2(_3652_),
    .C(_3526_),
    .ZN(_3661_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _8568_ (.A1(_3379_),
    .A2(_3645_),
    .B1(_3660_),
    .B2(_3661_),
    .C(_3373_),
    .ZN(_3662_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _8569_ (.A1(_2969_),
    .A2(_3621_),
    .B(_3662_),
    .C(_3592_),
    .ZN(_0218_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _8570_ (.A1(_2968_),
    .A2(_3644_),
    .ZN(_3663_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _8571_ (.A1(_0996_),
    .A2(_3663_),
    .Z(_3664_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _8572_ (.I(_3664_),
    .Z(_3665_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _8573_ (.A1(_0989_),
    .A2(_3648_),
    .ZN(_3666_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _8574_ (.A1(_0996_),
    .A2(_3666_),
    .Z(_3667_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _8575_ (.A1(_2950_),
    .A2(_3610_),
    .B(_2369_),
    .ZN(_3668_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_4 _8576_ (.A1(_2998_),
    .A2(_2538_),
    .A3(_3021_),
    .A4(_3609_),
    .ZN(_3669_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _8577_ (.A1(_3668_),
    .A2(_3669_),
    .ZN(_3670_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _8578_ (.A1(_3392_),
    .A2(_3665_),
    .ZN(_3671_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _8579_ (.A1(_3459_),
    .A2(_3667_),
    .B1(_3670_),
    .B2(_3504_),
    .C(_3671_),
    .ZN(_3672_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _8580_ (.I0(_0996_),
    .I1(_3006_),
    .S(_0837_),
    .Z(_3673_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _8581_ (.A1(_3533_),
    .A2(_3673_),
    .ZN(_3674_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _8582_ (.A1(_2368_),
    .A2(_2385_),
    .B(_3441_),
    .ZN(_3675_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _8583_ (.A1(_2481_),
    .A2(_2354_),
    .ZN(_3676_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _8584_ (.A1(_2495_),
    .A2(_3665_),
    .B1(_3675_),
    .B2(_1277_),
    .C(_3676_),
    .ZN(_3677_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _8585_ (.A1(_3256_),
    .A2(_3664_),
    .B1(_3673_),
    .B2(_2524_),
    .C(_2927_),
    .ZN(_3678_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _8586_ (.A1(_3674_),
    .A2(_3677_),
    .B(_3678_),
    .ZN(_3679_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _8587_ (.A1(_3153_),
    .A2(_3672_),
    .B(_3679_),
    .ZN(_3680_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _8588_ (.A1(_0533_),
    .A2(_3327_),
    .B1(_3317_),
    .B2(_3665_),
    .ZN(_3681_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _8589_ (.A1(_3680_),
    .A2(_3681_),
    .B(_3526_),
    .ZN(_3682_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _8590_ (.A1(_3292_),
    .A2(_3665_),
    .B(_3682_),
    .C(_3331_),
    .ZN(_3683_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _8591_ (.A1(_2995_),
    .A2(_3621_),
    .B(_3683_),
    .C(_3592_),
    .ZN(_0219_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _8592_ (.A1(\as2650.pc[11] ),
    .A2(_3663_),
    .ZN(_3684_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _8593_ (.A1(_3035_),
    .A2(_3684_),
    .Z(_3685_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _8594_ (.I(_3685_),
    .Z(_3686_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _8595_ (.A1(_0995_),
    .A2(_0988_),
    .A3(_3648_),
    .ZN(_3687_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _8596_ (.A1(_1003_),
    .A2(_3687_),
    .Z(_3688_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _8597_ (.A1(_3020_),
    .A2(_3669_),
    .Z(_3689_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _8598_ (.A1(_3394_),
    .A2(_3688_),
    .B1(_3689_),
    .B2(_3471_),
    .ZN(_3690_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _8599_ (.I0(_1002_),
    .I1(_3017_),
    .S(_1599_),
    .Z(_3691_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _8600_ (.A1(_2353_),
    .A2(_3691_),
    .ZN(_3692_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _8601_ (.A1(_2372_),
    .A2(_2776_),
    .B(_3470_),
    .ZN(_3693_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _8602_ (.A1(_3082_),
    .A2(_3686_),
    .B1(_3693_),
    .B2(_1276_),
    .C(_3676_),
    .ZN(_3694_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _8603_ (.A1(_3256_),
    .A2(_3685_),
    .B1(_3691_),
    .B2(_2523_),
    .C(_2855_),
    .ZN(_3695_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _8604_ (.A1(_3692_),
    .A2(_3694_),
    .B(_3695_),
    .ZN(_3696_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _8605_ (.A1(_3194_),
    .A2(_3690_),
    .B(_3696_),
    .ZN(_3697_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _8606_ (.A1(_3046_),
    .A2(_3697_),
    .ZN(_3698_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _8607_ (.A1(_3458_),
    .A2(_3686_),
    .B(_3698_),
    .ZN(_3699_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _8608_ (.A1(_0632_),
    .A2(_1499_),
    .B(_3699_),
    .ZN(_3700_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _8609_ (.A1(_3210_),
    .A2(_3686_),
    .B(_3700_),
    .ZN(_3701_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _8610_ (.A1(_3492_),
    .A2(_3686_),
    .B(_3331_),
    .ZN(_3702_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _8611_ (.A1(_3035_),
    .A2(_3374_),
    .B1(_3701_),
    .B2(_3702_),
    .C(_2415_),
    .ZN(_0220_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _8612_ (.I(_2415_),
    .Z(_3703_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _8613_ (.A1(_1002_),
    .A2(_0995_),
    .A3(_3663_),
    .ZN(_3704_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _8614_ (.A1(\as2650.pc[13] ),
    .A2(_3704_),
    .ZN(_3705_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _8615_ (.I(_3705_),
    .Z(_3706_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _8616_ (.A1(_3035_),
    .A2(_3687_),
    .ZN(_3707_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _8617_ (.A1(\as2650.pc[13] ),
    .A2(_3707_),
    .Z(_3708_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _8618_ (.I0(_3708_),
    .I1(_3705_),
    .S(_3353_),
    .Z(_3709_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _8619_ (.A1(_1251_),
    .A2(_3709_),
    .ZN(_3710_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _8620_ (.A1(_2996_),
    .A2(_3705_),
    .ZN(_3711_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _8621_ (.A1(_1008_),
    .A2(_1544_),
    .Z(_3712_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _8622_ (.A1(_4265_),
    .A2(_3345_),
    .B1(_2353_),
    .B2(_3712_),
    .C(_3048_),
    .ZN(_3713_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _8623_ (.A1(_3710_),
    .A2(_3711_),
    .A3(_3713_),
    .ZN(_3714_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _8624_ (.A1(_3093_),
    .A2(_3714_),
    .ZN(_3715_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _8625_ (.A1(_2372_),
    .A2(_3669_),
    .B(_3500_),
    .C(_2382_),
    .ZN(_3716_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _8626_ (.A1(_2926_),
    .A2(_3706_),
    .B(_3716_),
    .C(_3598_),
    .ZN(_3717_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _8627_ (.A1(_3257_),
    .A2(_3706_),
    .B1(_3712_),
    .B2(_2549_),
    .C(_2856_),
    .ZN(_3718_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _8628_ (.A1(_3715_),
    .A2(_3717_),
    .B(_3718_),
    .ZN(_3719_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _8629_ (.A1(_0709_),
    .A2(_3481_),
    .B1(_3426_),
    .B2(_3706_),
    .C(_3719_),
    .ZN(_3720_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _8630_ (.A1(_3329_),
    .A2(_3706_),
    .ZN(_3721_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _8631_ (.A1(_3379_),
    .A2(_3720_),
    .B(_3721_),
    .C(_3420_),
    .ZN(_3722_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _8632_ (.A1(_1008_),
    .A2(_3377_),
    .B(_3722_),
    .ZN(_3723_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _8633_ (.A1(_3703_),
    .A2(_3723_),
    .ZN(_0221_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _8634_ (.I(\as2650.pc[14] ),
    .ZN(_3724_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _8635_ (.A1(\as2650.pc[13] ),
    .A2(_1002_),
    .A3(_0995_),
    .A4(_3663_),
    .ZN(_3725_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _8636_ (.A1(_3724_),
    .A2(_3725_),
    .Z(_3726_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _8637_ (.I(_3726_),
    .Z(_3727_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _8638_ (.A1(_4264_),
    .A2(_3158_),
    .B(_3625_),
    .ZN(_3728_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _8639_ (.A1(_1008_),
    .A2(_3707_),
    .ZN(_3729_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _8640_ (.A1(\as2650.pc[14] ),
    .A2(_3729_),
    .Z(_3730_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _8641_ (.I(_3081_),
    .ZN(_3731_));
 gf180mcu_fd_sc_mcu7t5v0__aoi222_1 _8642_ (.A1(_4264_),
    .A2(_2410_),
    .B1(_2494_),
    .B2(_3726_),
    .C1(_3731_),
    .C2(\as2650.pc[14] ),
    .ZN(_3732_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _8643_ (.A1(_3430_),
    .A2(_3730_),
    .B1(_3732_),
    .B2(_2482_),
    .ZN(_3733_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _8644_ (.A1(_3393_),
    .A2(_3727_),
    .B1(_3733_),
    .B2(_3598_),
    .ZN(_3734_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _8645_ (.A1(_3728_),
    .A2(_3734_),
    .B(_3293_),
    .ZN(_3735_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _8646_ (.A1(_2634_),
    .A2(_3727_),
    .ZN(_3736_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _8647_ (.A1(_3724_),
    .A2(_3148_),
    .B(_3736_),
    .C(_3194_),
    .ZN(_3737_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _8648_ (.A1(_3214_),
    .A2(_3735_),
    .A3(_3737_),
    .ZN(_3738_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _8649_ (.A1(_0781_),
    .A2(_3327_),
    .B1(_2388_),
    .B2(_3727_),
    .ZN(_3739_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _8650_ (.A1(_3738_),
    .A2(_3739_),
    .B(_3526_),
    .ZN(_3740_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _8651_ (.A1(_3292_),
    .A2(_3727_),
    .B(_3740_),
    .C(_3373_),
    .ZN(_3741_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _8652_ (.I(_2577_),
    .Z(_3742_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _8653_ (.A1(_3724_),
    .A2(_3621_),
    .B(_3741_),
    .C(_3742_),
    .ZN(_0222_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _8654_ (.A1(_1453_),
    .A2(_2420_),
    .ZN(_3743_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _8655_ (.A1(_1329_),
    .A2(_2472_),
    .B(_3265_),
    .ZN(_3744_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_2 _8656_ (.A1(_2755_),
    .A2(_0600_),
    .B1(_3744_),
    .B2(_3175_),
    .C(_4260_),
    .ZN(_3745_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _8657_ (.A1(_3743_),
    .A2(_3745_),
    .B(_1516_),
    .ZN(_3746_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _8658_ (.A1(_4160_),
    .A2(_3265_),
    .A3(_1288_),
    .ZN(_3747_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _8659_ (.A1(_2927_),
    .A2(_3747_),
    .B(_0971_),
    .ZN(_3748_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _8660_ (.A1(_4419_),
    .A2(_1046_),
    .B(_4395_),
    .ZN(_3749_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_2 _8661_ (.A1(_1463_),
    .A2(_3748_),
    .B1(_3749_),
    .B2(_3265_),
    .ZN(_3750_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _8662_ (.A1(_1328_),
    .A2(_1338_),
    .B(_1496_),
    .C(_2448_),
    .ZN(_3751_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_1 _8663_ (.A1(_4242_),
    .A2(_2469_),
    .A3(_1491_),
    .B(_3751_),
    .ZN(_3752_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _8664_ (.I(_3752_),
    .ZN(_3753_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_2 _8665_ (.A1(_1939_),
    .A2(_0871_),
    .A3(_1352_),
    .A4(_1487_),
    .ZN(_3754_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_2 _8666_ (.A1(_1333_),
    .A2(_1474_),
    .A3(_3753_),
    .A4(_3754_),
    .ZN(_3755_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_2 _8667_ (.A1(_1318_),
    .A2(_1476_),
    .A3(_1478_),
    .A4(_1484_),
    .ZN(_3756_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_4 _8668_ (.A1(_3746_),
    .A2(_3750_),
    .A3(_3755_),
    .A4(_3756_),
    .ZN(_3757_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _8669_ (.I(_3757_),
    .Z(_3758_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _8670_ (.A1(_2598_),
    .A2(_4361_),
    .ZN(_3759_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _8671_ (.A1(_2477_),
    .A2(_4353_),
    .B(_3759_),
    .ZN(_3760_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _8672_ (.A1(_3143_),
    .A2(_1100_),
    .B(_3080_),
    .ZN(_3761_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_1 _8673_ (.A1(_3219_),
    .A2(_4344_),
    .B1(_3183_),
    .B2(_3760_),
    .C(_3761_),
    .ZN(_3762_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _8674_ (.I(_3757_),
    .Z(_3763_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _8675_ (.A1(_4398_),
    .A2(_2632_),
    .ZN(_3764_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _8676_ (.I(_4394_),
    .Z(_3765_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _8677_ (.I(_3765_),
    .Z(_3766_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _8678_ (.I(_1535_),
    .Z(_3767_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _8679_ (.A1(_0618_),
    .A2(_3326_),
    .ZN(_3768_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _8680_ (.I(_1235_),
    .Z(_3769_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _8681_ (.A1(_4428_),
    .A2(_4137_),
    .ZN(_3770_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_2 _8682_ (.A1(_0550_),
    .A2(_3770_),
    .A3(_0340_),
    .ZN(_3771_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _8683_ (.I(_3771_),
    .Z(_3772_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _8684_ (.I(_3771_),
    .Z(_3773_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _8685_ (.A1(_1589_),
    .A2(_3773_),
    .ZN(_3774_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _8686_ (.A1(_4316_),
    .A2(_3772_),
    .B(_3774_),
    .ZN(_3775_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _8687_ (.A1(_1736_),
    .A2(_3769_),
    .B1(_4435_),
    .B2(_3775_),
    .ZN(_3776_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _8688_ (.I(_4219_),
    .Z(_3777_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _8689_ (.A1(_3768_),
    .A2(_3776_),
    .B(_3777_),
    .ZN(_3778_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _8690_ (.A1(_1624_),
    .A2(_4377_),
    .B(_3778_),
    .C(_1535_),
    .ZN(_3779_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _8691_ (.I(_4394_),
    .Z(_3780_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _8692_ (.A1(_3767_),
    .A2(_1383_),
    .B(_3779_),
    .C(_3780_),
    .ZN(_3781_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _8693_ (.A1(_1691_),
    .A2(_3766_),
    .B(_2629_),
    .C(_3781_),
    .ZN(_3782_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _8694_ (.A1(_3762_),
    .A2(_3763_),
    .A3(_3764_),
    .A4(_3782_),
    .ZN(_3783_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _8695_ (.A1(_4441_),
    .A2(_3758_),
    .B(_3783_),
    .ZN(_3784_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _8696_ (.A1(_3703_),
    .A2(_3784_),
    .ZN(_0223_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _8697_ (.I(_2337_),
    .Z(_3785_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _8698_ (.I0(_4513_),
    .I1(_0292_),
    .S(_3785_),
    .Z(_3786_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _8699_ (.A1(_3143_),
    .A2(_1383_),
    .B(_3080_),
    .ZN(_3787_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_1 _8700_ (.A1(_3219_),
    .A2(_0321_),
    .B1(_3183_),
    .B2(_3786_),
    .C(_3787_),
    .ZN(_3788_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _8701_ (.A1(_1552_),
    .A2(_1541_),
    .B(_3170_),
    .ZN(_3789_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _8702_ (.I(_4227_),
    .Z(_3790_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _8703_ (.A1(_0619_),
    .A2(_3368_),
    .ZN(_3791_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _8704_ (.I(_2423_),
    .Z(_3792_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _8705_ (.I(_3792_),
    .Z(_3793_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _8706_ (.A1(\as2650.psl[1] ),
    .A2(_3792_),
    .ZN(_3794_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _8707_ (.A1(_4458_),
    .A2(_3793_),
    .B(_3794_),
    .ZN(_3795_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_1 _8708_ (.A1(_1733_),
    .A2(_3769_),
    .B1(_4435_),
    .B2(_3795_),
    .C(_3777_),
    .ZN(_3796_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _8709_ (.A1(_1519_),
    .A2(_4514_),
    .B(_1480_),
    .ZN(_3797_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _8710_ (.A1(_3791_),
    .A2(_3796_),
    .B(_3797_),
    .ZN(_3798_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _8711_ (.A1(_3790_),
    .A2(_0400_),
    .B(_3798_),
    .C(_3765_),
    .ZN(_3799_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _8712_ (.A1(_3199_),
    .A2(_4535_),
    .B1(_3789_),
    .B2(_3799_),
    .ZN(_3800_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _8713_ (.A1(_3088_),
    .A2(_3800_),
    .ZN(_3801_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _8714_ (.A1(_3763_),
    .A2(_3788_),
    .A3(_3801_),
    .ZN(_3802_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _8715_ (.A1(_1382_),
    .A2(_3758_),
    .B(_3802_),
    .ZN(_3803_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _8716_ (.A1(_3703_),
    .A2(_3803_),
    .ZN(_0224_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _8717_ (.I(_2337_),
    .Z(_3804_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _8718_ (.A1(_3785_),
    .A2(_0358_),
    .ZN(_3805_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _8719_ (.A1(_3804_),
    .A2(_2592_),
    .B(_3805_),
    .ZN(_3806_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _8720_ (.A1(_3143_),
    .A2(_4527_),
    .B(_3080_),
    .ZN(_3807_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_1 _8721_ (.A1(_3219_),
    .A2(_0422_),
    .B1(_3183_),
    .B2(_3806_),
    .C(_3807_),
    .ZN(_3808_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _8722_ (.A1(_0378_),
    .A2(_2632_),
    .ZN(_3809_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _8723_ (.I(_1623_),
    .Z(_3810_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _8724_ (.A1(_0618_),
    .A2(_3390_),
    .ZN(_3811_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _8725_ (.I(\as2650.overflow ),
    .ZN(_3812_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _8726_ (.A1(_0849_),
    .A2(_3773_),
    .ZN(_3813_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _8727_ (.A1(_3812_),
    .A2(_3772_),
    .B(_3813_),
    .ZN(_3814_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_1 _8728_ (.A1(_3769_),
    .A2(_1749_),
    .B1(_3814_),
    .B2(_4435_),
    .C(_1623_),
    .ZN(_3815_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _8729_ (.A1(_3810_),
    .A2(_4388_),
    .B1(_3811_),
    .B2(_3815_),
    .ZN(_3816_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _8730_ (.A1(_3790_),
    .A2(_3816_),
    .ZN(_3817_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _8731_ (.A1(_3767_),
    .A2(_1393_),
    .B(_3817_),
    .C(_3765_),
    .ZN(_3818_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _8732_ (.A1(_1699_),
    .A2(_3766_),
    .B(_2629_),
    .C(_3818_),
    .ZN(_3819_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _8733_ (.A1(_3763_),
    .A2(_3808_),
    .A3(_3809_),
    .A4(_3819_),
    .ZN(_3820_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _8734_ (.A1(_0917_),
    .A2(_3758_),
    .B(_3820_),
    .ZN(_3821_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _8735_ (.A1(_3703_),
    .A2(_3821_),
    .ZN(_0225_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _8736_ (.A1(_2338_),
    .A2(_0491_),
    .ZN(_3822_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _8737_ (.A1(_3785_),
    .A2(_0485_),
    .B(_3822_),
    .C(_2756_),
    .ZN(_3823_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _8738_ (.A1(_2756_),
    .A2(_0476_),
    .B(_3823_),
    .C(_3126_),
    .ZN(_3824_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _8739_ (.A1(_3144_),
    .A2(_1393_),
    .B(_3824_),
    .C(_3088_),
    .ZN(_3825_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _8740_ (.A1(_0618_),
    .A2(_3451_),
    .ZN(_3826_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _8741_ (.I(_4365_),
    .ZN(_3827_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _8742_ (.A1(\as2650.psu[3] ),
    .A2(_3771_),
    .ZN(_3828_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _8743_ (.A1(_3827_),
    .A2(_3773_),
    .B(_3828_),
    .ZN(_3829_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _8744_ (.A1(_1235_),
    .A2(_1764_),
    .B1(_3829_),
    .B2(_4434_),
    .ZN(_3830_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _8745_ (.A1(_3826_),
    .A2(_3830_),
    .B(_3777_),
    .ZN(_3831_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _8746_ (.A1(_3810_),
    .A2(_0400_),
    .B(_3831_),
    .C(_1535_),
    .ZN(_3832_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _8747_ (.A1(_3790_),
    .A2(_0694_),
    .B(_3832_),
    .C(_3765_),
    .ZN(_3833_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _8748_ (.A1(_1556_),
    .A2(_3780_),
    .B(_2629_),
    .C(_3833_),
    .ZN(_3834_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _8749_ (.A1(_0512_),
    .A2(_2753_),
    .B(_3757_),
    .C(_3834_),
    .ZN(_3835_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _8750_ (.A1(_0924_),
    .A2(_3758_),
    .B1(_3825_),
    .B2(_3835_),
    .ZN(_3836_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _8751_ (.A1(_3189_),
    .A2(_3836_),
    .ZN(_0226_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _8752_ (.I(_3763_),
    .Z(_3837_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _8753_ (.I(_2386_),
    .Z(_3838_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _8754_ (.A1(_3804_),
    .A2(_0614_),
    .Z(_3839_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _8755_ (.A1(_2477_),
    .A2(_0578_),
    .B(_3839_),
    .ZN(_3840_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _8756_ (.A1(_1572_),
    .A2(_0566_),
    .B(_1518_),
    .ZN(_3841_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_1 _8757_ (.A1(_3838_),
    .A2(_0570_),
    .B1(_3184_),
    .B2(_3840_),
    .C(_3841_),
    .ZN(_3842_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _8758_ (.A1(_0619_),
    .A2(_3488_),
    .ZN(_3843_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _8759_ (.I(_1235_),
    .Z(_3844_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _8760_ (.A1(\as2650.psu[4] ),
    .A2(_3772_),
    .ZN(_3845_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _8761_ (.A1(_1033_),
    .A2(_3772_),
    .B(_3845_),
    .ZN(_3846_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _8762_ (.I(_4434_),
    .Z(_3847_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_1 _8763_ (.A1(_3844_),
    .A2(_2027_),
    .B1(_3846_),
    .B2(_3847_),
    .C(_3810_),
    .ZN(_3848_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _8764_ (.A1(_1520_),
    .A2(_0372_),
    .ZN(_3849_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _8765_ (.A1(_3843_),
    .A2(_3848_),
    .B(_3849_),
    .C(_3767_),
    .ZN(_3850_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _8766_ (.I(_1628_),
    .Z(_3851_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _8767_ (.A1(_3851_),
    .A2(_0593_),
    .B(_1541_),
    .ZN(_3852_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _8768_ (.A1(_1558_),
    .A2(_1547_),
    .B1(_3850_),
    .B2(_3852_),
    .C(_1513_),
    .ZN(_3853_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _8769_ (.A1(_0603_),
    .A2(_2633_),
    .B(_3853_),
    .ZN(_3854_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _8770_ (.A1(_3842_),
    .A2(_3854_),
    .ZN(_3855_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _8771_ (.I(_3757_),
    .Z(_3856_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _8772_ (.A1(_0579_),
    .A2(_3856_),
    .B(_3245_),
    .ZN(_3857_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _8773_ (.A1(_3837_),
    .A2(_3855_),
    .B(_3857_),
    .ZN(_0227_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _8774_ (.A1(_2598_),
    .A2(_0698_),
    .Z(_3858_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _8775_ (.A1(_3804_),
    .A2(_0668_),
    .B(_3858_),
    .ZN(_3859_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _8776_ (.A1(_2399_),
    .A2(_0639_),
    .B(_2514_),
    .ZN(_3860_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_1 _8777_ (.A1(_3838_),
    .A2(_0662_),
    .B1(_3184_),
    .B2(_3859_),
    .C(_3860_),
    .ZN(_3861_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _8778_ (.A1(_3810_),
    .A2(_0694_),
    .ZN(_3862_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _8779_ (.A1(\as2650.psl[5] ),
    .A2(_3792_),
    .ZN(_3863_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _8780_ (.A1(_1226_),
    .A2(_3793_),
    .B(_3863_),
    .ZN(_3864_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_1 _8781_ (.A1(_3769_),
    .A2(_1812_),
    .B1(_3864_),
    .B2(_3847_),
    .C(_1623_),
    .ZN(_3865_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _8782_ (.A1(_0341_),
    .A2(_3525_),
    .B(_3865_),
    .ZN(_3866_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _8783_ (.A1(_3862_),
    .A2(_3866_),
    .B(_3790_),
    .ZN(_3867_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _8784_ (.A1(_1628_),
    .A2(_1537_),
    .ZN(_3868_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _8785_ (.A1(_3780_),
    .A2(_3867_),
    .A3(_3868_),
    .ZN(_3869_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _8786_ (.A1(_1292_),
    .A2(_3766_),
    .B(_3869_),
    .ZN(_3870_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _8787_ (.A1(_0690_),
    .A2(_2633_),
    .B1(_3870_),
    .B2(_2630_),
    .ZN(_3871_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _8788_ (.A1(_3861_),
    .A2(_3871_),
    .ZN(_3872_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _8789_ (.A1(_0711_),
    .A2(_3856_),
    .B(_3245_),
    .ZN(_3873_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _8790_ (.A1(_3837_),
    .A2(_3872_),
    .B(_3873_),
    .ZN(_0228_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _8791_ (.A1(_2565_),
    .A2(_0771_),
    .Z(_3874_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _8792_ (.A1(_3804_),
    .A2(_0749_),
    .B(_3874_),
    .ZN(_3875_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _8793_ (.A1(_2635_),
    .A2(_1537_),
    .B(_1450_),
    .ZN(_3876_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_1 _8794_ (.A1(_3838_),
    .A2(_0740_),
    .B1(_3184_),
    .B2(_3875_),
    .C(_3876_),
    .ZN(_3877_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _8795_ (.I0(net27),
    .I1(_1525_),
    .S(_3792_),
    .Z(_3878_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_1 _8796_ (.A1(_3844_),
    .A2(_2084_),
    .B1(_3878_),
    .B2(_3847_),
    .C(_3777_),
    .ZN(_3879_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _8797_ (.A1(_0342_),
    .A2(_3557_),
    .B(_3879_),
    .ZN(_3880_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _8798_ (.A1(_1627_),
    .A2(_0639_),
    .B(_3880_),
    .C(_3851_),
    .ZN(_3881_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _8799_ (.A1(_3767_),
    .A2(_0818_),
    .B(_3780_),
    .ZN(_3882_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_1 _8800_ (.A1(_1588_),
    .A2(_3766_),
    .B1(_3881_),
    .B2(_3882_),
    .C(_2630_),
    .ZN(_3883_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _8801_ (.A1(_2458_),
    .A2(_2753_),
    .B(_3877_),
    .C(_3883_),
    .ZN(_3884_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _8802_ (.A1(_0944_),
    .A2(_3856_),
    .B(_3245_),
    .ZN(_3885_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _8803_ (.A1(_3837_),
    .A2(_3884_),
    .B(_3885_),
    .ZN(_0229_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _8804_ (.A1(_2338_),
    .A2(_0830_),
    .ZN(_3886_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _8805_ (.A1(_3785_),
    .A2(_0828_),
    .B(_3182_),
    .C(_3886_),
    .ZN(_3887_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _8806_ (.A1(_2635_),
    .A2(_0818_),
    .B(_3887_),
    .C(_2514_),
    .ZN(_3888_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _8807_ (.A1(_3838_),
    .A2(_1212_),
    .B(_3888_),
    .ZN(_3889_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _8808_ (.A1(_0620_),
    .A2(_3588_),
    .ZN(_3890_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _8809_ (.A1(_1611_),
    .A2(_3793_),
    .ZN(_3891_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _8810_ (.A1(_3262_),
    .A2(_3793_),
    .B(_3891_),
    .ZN(_3892_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_1 _8811_ (.A1(_2109_),
    .A2(_3844_),
    .B1(_3847_),
    .B2(_3892_),
    .C(_1624_),
    .ZN(_3893_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _8812_ (.A1(_3890_),
    .A2(_3893_),
    .B(_1629_),
    .ZN(_3894_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _8813_ (.A1(_1577_),
    .A2(_3894_),
    .ZN(_3895_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _8814_ (.A1(_2630_),
    .A2(_1548_),
    .A3(_3895_),
    .ZN(_3896_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _8815_ (.A1(_0834_),
    .A2(_2753_),
    .B(_3889_),
    .C(_3896_),
    .ZN(_3897_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _8816_ (.A1(_1411_),
    .A2(_3856_),
    .B(_1634_),
    .ZN(_3898_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _8817_ (.A1(_3837_),
    .A2(_3897_),
    .B(_3898_),
    .ZN(_0230_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _8818_ (.A1(_0957_),
    .A2(_0427_),
    .ZN(_3899_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _8819_ (.A1(_2208_),
    .A2(_3899_),
    .ZN(_3900_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _8820_ (.I(_3900_),
    .Z(_3901_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _8821_ (.I(_3901_),
    .Z(_3902_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _8822_ (.A1(_0958_),
    .A2(_2212_),
    .ZN(_3903_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _8823_ (.I(_3903_),
    .Z(_3904_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _8824_ (.A1(_2223_),
    .A2(_0626_),
    .A3(_0901_),
    .ZN(_3905_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _8825_ (.I(_3905_),
    .Z(_3906_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _8826_ (.A1(_2146_),
    .A2(_3904_),
    .B1(_3906_),
    .B2(\as2650.stack[6][0] ),
    .C(_3901_),
    .ZN(_3907_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _8827_ (.A1(_0848_),
    .A2(_3902_),
    .B(_3907_),
    .ZN(_0231_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _8828_ (.I(_3903_),
    .Z(_3908_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _8829_ (.I(_3905_),
    .Z(_3909_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _8830_ (.I(_3900_),
    .Z(_3910_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _8831_ (.A1(_2285_),
    .A2(_3908_),
    .B1(_3909_),
    .B2(\as2650.stack[6][1] ),
    .C(_3910_),
    .ZN(_3911_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _8832_ (.A1(_2223_),
    .A2(_0624_),
    .A3(_0968_),
    .ZN(_3912_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _8833_ (.A1(_2290_),
    .A2(_3912_),
    .ZN(_3913_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _8834_ (.A1(_3911_),
    .A2(_3913_),
    .ZN(_0232_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _8835_ (.A1(_2258_),
    .A2(_3908_),
    .B1(_3909_),
    .B2(\as2650.stack[6][2] ),
    .C(_3910_),
    .ZN(_3914_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _8836_ (.A1(_2294_),
    .A2(_3912_),
    .ZN(_3915_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _8837_ (.A1(_3914_),
    .A2(_3915_),
    .ZN(_0233_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _8838_ (.A1(_2296_),
    .A2(_3908_),
    .B1(_3909_),
    .B2(\as2650.stack[6][3] ),
    .C(_3910_),
    .ZN(_3916_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _8839_ (.A1(_2298_),
    .A2(_3912_),
    .ZN(_3917_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _8840_ (.A1(_3916_),
    .A2(_3917_),
    .ZN(_0234_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _8841_ (.A1(_2300_),
    .A2(_3904_),
    .B1(_3906_),
    .B2(\as2650.stack[6][4] ),
    .C(_3901_),
    .ZN(_3918_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _8842_ (.A1(_0932_),
    .A2(_3902_),
    .B(_3918_),
    .ZN(_0235_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _8843_ (.A1(_2302_),
    .A2(_3904_),
    .B1(_3906_),
    .B2(\as2650.stack[6][5] ),
    .C(_3901_),
    .ZN(_3919_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _8844_ (.A1(_0938_),
    .A2(_3902_),
    .B(_3919_),
    .ZN(_0236_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _8845_ (.A1(_2265_),
    .A2(_3904_),
    .B1(_3906_),
    .B2(\as2650.stack[6][6] ),
    .C(_3910_),
    .ZN(_3920_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _8846_ (.A1(_2199_),
    .A2(_3902_),
    .B(_3920_),
    .ZN(_0237_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _8847_ (.A1(_2305_),
    .A2(_3908_),
    .B1(_3909_),
    .B2(\as2650.stack[6][7] ),
    .C(_3900_),
    .ZN(_3921_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _8848_ (.A1(_2307_),
    .A2(_3912_),
    .ZN(_3922_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _8849_ (.A1(_3921_),
    .A2(_3922_),
    .ZN(_0238_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _8850_ (.A1(_0857_),
    .A2(_2314_),
    .Z(_3923_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _8851_ (.I(_3923_),
    .Z(_3924_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _8852_ (.I(_3924_),
    .Z(_3925_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _8853_ (.A1(_2212_),
    .A2(_3899_),
    .ZN(_3926_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _8854_ (.I(_3926_),
    .Z(_3927_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _8855_ (.A1(_2148_),
    .A2(_0624_),
    .A3(_0901_),
    .ZN(_3928_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _8856_ (.I(_3928_),
    .Z(_3929_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _8857_ (.A1(_2146_),
    .A2(_3927_),
    .B1(_3929_),
    .B2(\as2650.stack[7][0] ),
    .C(_3924_),
    .ZN(_3930_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _8858_ (.A1(_0848_),
    .A2(_3925_),
    .B(_3930_),
    .ZN(_0239_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _8859_ (.I(_3926_),
    .Z(_3931_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _8860_ (.I(_3928_),
    .Z(_3932_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _8861_ (.I(_3923_),
    .Z(_3933_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _8862_ (.A1(_2285_),
    .A2(_3931_),
    .B1(_3932_),
    .B2(\as2650.stack[7][1] ),
    .C(_3933_),
    .ZN(_3934_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _8863_ (.A1(_0968_),
    .A2(_2314_),
    .ZN(_3935_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _8864_ (.A1(_2290_),
    .A2(_3935_),
    .ZN(_3936_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _8865_ (.A1(_3934_),
    .A2(_3936_),
    .ZN(_0240_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _8866_ (.A1(_0921_),
    .A2(_3931_),
    .B1(_3932_),
    .B2(\as2650.stack[7][2] ),
    .C(_3933_),
    .ZN(_3937_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _8867_ (.A1(_2294_),
    .A2(_3935_),
    .ZN(_3938_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _8868_ (.A1(_3937_),
    .A2(_3938_),
    .ZN(_0241_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _8869_ (.A1(_2296_),
    .A2(_3931_),
    .B1(_3932_),
    .B2(\as2650.stack[7][3] ),
    .C(_3933_),
    .ZN(_3939_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _8870_ (.A1(_2298_),
    .A2(_3935_),
    .ZN(_3940_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _8871_ (.A1(_3939_),
    .A2(_3940_),
    .ZN(_0242_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _8872_ (.A1(_2300_),
    .A2(_3927_),
    .B1(_3929_),
    .B2(\as2650.stack[7][4] ),
    .C(_3924_),
    .ZN(_3941_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _8873_ (.A1(_0932_),
    .A2(_3925_),
    .B(_3941_),
    .ZN(_0243_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _8874_ (.A1(_2302_),
    .A2(_3927_),
    .B1(_3929_),
    .B2(\as2650.stack[7][5] ),
    .C(_3924_),
    .ZN(_3942_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _8875_ (.A1(_0938_),
    .A2(_3925_),
    .B(_3942_),
    .ZN(_0244_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _8876_ (.A1(_0948_),
    .A2(_3927_),
    .B1(_3929_),
    .B2(\as2650.stack[7][6] ),
    .C(_3933_),
    .ZN(_3943_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _8877_ (.A1(_2199_),
    .A2(_3925_),
    .B(_3943_),
    .ZN(_0245_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _8878_ (.A1(_2305_),
    .A2(_3931_),
    .B1(_3932_),
    .B2(\as2650.stack[7][7] ),
    .C(_3923_),
    .ZN(_3944_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _8879_ (.A1(_2307_),
    .A2(_3935_),
    .ZN(_3945_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _8880_ (.A1(_3944_),
    .A2(_3945_),
    .ZN(_0246_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _8881_ (.A1(_1019_),
    .A2(_3899_),
    .ZN(_3946_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _8882_ (.I(_3946_),
    .Z(_3947_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _8883_ (.I(_3947_),
    .Z(_3948_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _8884_ (.I(_3947_),
    .Z(_3949_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _8885_ (.A1(\as2650.stack[7][8] ),
    .A2(_3949_),
    .ZN(_3950_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _8886_ (.A1(_1653_),
    .A2(_3948_),
    .B(_3950_),
    .ZN(_0247_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _8887_ (.I(_3946_),
    .Z(_3951_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _8888_ (.A1(\as2650.stack[7][9] ),
    .A2(_3951_),
    .ZN(_3952_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _8889_ (.A1(_1663_),
    .A2(_3948_),
    .B(_3952_),
    .ZN(_0248_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _8890_ (.A1(\as2650.stack[7][10] ),
    .A2(_3951_),
    .ZN(_3953_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _8891_ (.A1(_1666_),
    .A2(_3948_),
    .B(_3953_),
    .ZN(_0249_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _8892_ (.A1(\as2650.stack[7][11] ),
    .A2(_3951_),
    .ZN(_3954_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _8893_ (.A1(_1668_),
    .A2(_3948_),
    .B(_3954_),
    .ZN(_0250_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _8894_ (.A1(\as2650.stack[7][12] ),
    .A2(_3951_),
    .ZN(_3955_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _8895_ (.A1(_1670_),
    .A2(_3949_),
    .B(_3955_),
    .ZN(_0251_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _8896_ (.A1(\as2650.stack[7][13] ),
    .A2(_3947_),
    .ZN(_3956_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _8897_ (.A1(_1672_),
    .A2(_3949_),
    .B(_3956_),
    .ZN(_0252_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _8898_ (.A1(\as2650.stack[7][14] ),
    .A2(_3947_),
    .ZN(_3957_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _8899_ (.A1(_1674_),
    .A2(_3949_),
    .B(_3957_),
    .ZN(_0253_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _8900_ (.A1(_1601_),
    .A2(_4272_),
    .ZN(_3958_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _8901_ (.I(_3958_),
    .ZN(_3959_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _8902_ (.A1(_4153_),
    .A2(_4491_),
    .ZN(_3960_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _8903_ (.I(_3960_),
    .Z(_3961_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _8904_ (.I(_3961_),
    .Z(_3962_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _8905_ (.A1(_1390_),
    .A2(_3960_),
    .A3(_3958_),
    .ZN(_3963_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _8906_ (.I(_3963_),
    .Z(_3964_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _8907_ (.A1(_3962_),
    .A2(_1724_),
    .B1(_3964_),
    .B2(\as2650.r123[1][0] ),
    .ZN(_3965_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _8908_ (.A1(_4414_),
    .A2(_3959_),
    .B(_3965_),
    .ZN(_0254_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _8909_ (.I(_3961_),
    .Z(_3966_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _8910_ (.I(_3963_),
    .Z(_3967_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _8911_ (.A1(_3966_),
    .A2(_1738_),
    .B1(_3967_),
    .B2(\as2650.r123[1][1] ),
    .ZN(_3968_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _8912_ (.I(_3958_),
    .Z(_3969_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _8913_ (.A1(_0323_),
    .A2(_3969_),
    .ZN(_3970_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _8914_ (.A1(_3968_),
    .A2(_3970_),
    .ZN(_0255_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _8915_ (.A1(_3966_),
    .A2(_1753_),
    .B1(_3967_),
    .B2(\as2650.r123[1][2] ),
    .ZN(_3971_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _8916_ (.A1(_0424_),
    .A2(_3969_),
    .ZN(_3972_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _8917_ (.A1(_3971_),
    .A2(_3972_),
    .ZN(_0256_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _8918_ (.A1(_3962_),
    .A2(_1772_),
    .B1(_3964_),
    .B2(\as2650.r123[1][3] ),
    .ZN(_3973_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _8919_ (.A1(_0523_),
    .A2(_3959_),
    .B(_3973_),
    .ZN(_0257_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _8920_ (.A1(_3962_),
    .A2(_1792_),
    .B1(_3964_),
    .B2(\as2650.r123[1][4] ),
    .ZN(_3974_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _8921_ (.A1(_0616_),
    .A2(_3969_),
    .ZN(_3975_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _8922_ (.A1(_3974_),
    .A2(_3975_),
    .ZN(_0258_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _8923_ (.A1(_0981_),
    .A2(_1939_),
    .ZN(_3976_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _8924_ (.A1(_3976_),
    .A2(_1823_),
    .ZN(_3977_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _8925_ (.A1(\as2650.r123[1][5] ),
    .A2(_3967_),
    .B(_3977_),
    .ZN(_3978_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _8926_ (.A1(_0703_),
    .A2(_3969_),
    .ZN(_3979_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _8927_ (.A1(_3978_),
    .A2(_3979_),
    .ZN(_0259_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _8928_ (.A1(_3976_),
    .A2(_1859_),
    .ZN(_3980_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _8929_ (.A1(\as2650.r123[1][6] ),
    .A2(_3967_),
    .B(_3980_),
    .ZN(_3981_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _8930_ (.A1(_0775_),
    .A2(_3958_),
    .ZN(_3982_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _8931_ (.A1(_3981_),
    .A2(_3982_),
    .ZN(_0260_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _8932_ (.A1(_3976_),
    .A2(_1898_),
    .ZN(_3983_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _8933_ (.A1(\as2650.r123[1][7] ),
    .A2(_3964_),
    .B(_3983_),
    .ZN(_3984_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _8934_ (.A1(_0846_),
    .A2(_3959_),
    .B(_3984_),
    .ZN(_0261_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _8935_ (.A1(_4272_),
    .A2(_1612_),
    .ZN(_3985_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _8936_ (.I(_3985_),
    .Z(_3986_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _8937_ (.I(_3986_),
    .ZN(_3987_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _8938_ (.A1(_1390_),
    .A2(_3961_),
    .A3(_3985_),
    .ZN(_3988_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _8939_ (.I(_3988_),
    .Z(_3989_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _8940_ (.A1(\as2650.r123[2][0] ),
    .A2(_3989_),
    .ZN(_3990_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _8941_ (.A1(_3966_),
    .A2(_1979_),
    .ZN(_3991_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _8942_ (.A1(_4414_),
    .A2(_3987_),
    .B(_3990_),
    .C(_3991_),
    .ZN(_0262_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _8943_ (.I(_3986_),
    .Z(_3992_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _8944_ (.I(_3988_),
    .Z(_3993_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _8945_ (.A1(_0323_),
    .A2(_3992_),
    .B1(_3993_),
    .B2(\as2650.r123[2][1] ),
    .ZN(_3994_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _8946_ (.I(_3961_),
    .Z(_3995_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _8947_ (.A1(_3995_),
    .A2(_2017_),
    .ZN(_3996_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _8948_ (.A1(_3994_),
    .A2(_3996_),
    .ZN(_0263_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _8949_ (.A1(_0424_),
    .A2(_3992_),
    .B1(_3993_),
    .B2(\as2650.r123[2][2] ),
    .ZN(_3997_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _8950_ (.A1(_3995_),
    .A2(_2048_),
    .ZN(_3998_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _8951_ (.A1(_3997_),
    .A2(_3998_),
    .ZN(_0264_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _8952_ (.A1(_0524_),
    .A2(_3992_),
    .B1(_3993_),
    .B2(\as2650.r123[2][3] ),
    .ZN(_3999_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _8953_ (.A1(_3995_),
    .A2(_2076_),
    .ZN(_4000_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _8954_ (.A1(_3999_),
    .A2(_4000_),
    .ZN(_0265_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _8955_ (.A1(_0616_),
    .A2(_3986_),
    .B1(_3989_),
    .B2(\as2650.r123[2][4] ),
    .ZN(_4001_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _8956_ (.A1(_3976_),
    .A2(_2100_),
    .B(_4001_),
    .ZN(_0266_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _8957_ (.A1(_0703_),
    .A2(_3992_),
    .B1(_3993_),
    .B2(\as2650.r123[2][5] ),
    .ZN(_4002_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _8958_ (.A1(_3995_),
    .A2(_2117_),
    .ZN(_4003_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _8959_ (.A1(_4002_),
    .A2(_4003_),
    .ZN(_0267_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _8960_ (.A1(_0775_),
    .A2(_3986_),
    .B1(_3989_),
    .B2(\as2650.r123[2][6] ),
    .ZN(_4004_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _8961_ (.A1(_3966_),
    .A2(_2129_),
    .ZN(_4005_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _8962_ (.A1(_4004_),
    .A2(_4005_),
    .ZN(_0268_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _8963_ (.A1(\as2650.r123[2][7] ),
    .A2(_3989_),
    .ZN(_4006_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_1 _8964_ (.A1(_2131_),
    .A2(_2132_),
    .A3(_2135_),
    .B(_3962_),
    .ZN(_4007_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _8965_ (.A1(_0846_),
    .A2(_3987_),
    .B(_4006_),
    .C(_4007_),
    .ZN(_0269_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _8966_ (.A1(_1556_),
    .A2(_1704_),
    .ZN(_4008_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _8967_ (.A1(_3191_),
    .A2(_1698_),
    .B(_4008_),
    .ZN(_0270_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _8968_ (.A1(_2373_),
    .A2(_1704_),
    .ZN(_4009_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _8969_ (.A1(_1570_),
    .A2(_1698_),
    .B(_4009_),
    .ZN(_0271_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _8970_ (.A1(_1555_),
    .A2(_2634_),
    .ZN(_4010_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_1 _8971_ (.A1(_3191_),
    .A2(_2509_),
    .A3(_3048_),
    .A4(_1309_),
    .ZN(_4011_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _8972_ (.A1(_2926_),
    .A2(_4011_),
    .ZN(_4012_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _8973_ (.A1(_2409_),
    .A2(_1481_),
    .ZN(_4013_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_1 _8974_ (.A1(_3045_),
    .A2(_1246_),
    .B1(_1265_),
    .B2(_4013_),
    .C(_3273_),
    .ZN(_4014_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _8975_ (.I(_4014_),
    .ZN(_4015_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _8976_ (.A1(_1482_),
    .A2(_3163_),
    .A3(_0875_),
    .ZN(_4016_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _8977_ (.A1(_1250_),
    .A2(_3773_),
    .ZN(_4017_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _8978_ (.A1(_4017_),
    .A2(_1467_),
    .ZN(_4018_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _8979_ (.A1(_1278_),
    .A2(_1242_),
    .B(_1716_),
    .C(_4018_),
    .ZN(_4019_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _8980_ (.A1(_2342_),
    .A2(_2400_),
    .A3(_4016_),
    .A4(_4019_),
    .ZN(_4020_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _8981_ (.A1(_3057_),
    .A2(_0897_),
    .B1(_2408_),
    .B2(_1272_),
    .ZN(_4021_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _8982_ (.A1(_1498_),
    .A2(_3236_),
    .B(_4021_),
    .ZN(_4022_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _8983_ (.A1(_3844_),
    .A2(_2449_),
    .A3(_1281_),
    .A4(_1357_),
    .ZN(_4023_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_2 _8984_ (.A1(_1046_),
    .A2(_4020_),
    .A3(_4022_),
    .A4(_4023_),
    .ZN(_4024_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_2 _8985_ (.A1(_3415_),
    .A2(_2438_),
    .B(_3084_),
    .C(_3275_),
    .ZN(_4025_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_2 _8986_ (.A1(_4012_),
    .A2(_4015_),
    .A3(_4024_),
    .A4(_4025_),
    .ZN(_4026_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _8987_ (.A1(_3336_),
    .A2(_4010_),
    .B(_4026_),
    .ZN(_4027_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _8988_ (.A1(_2634_),
    .A2(_3266_),
    .ZN(_4028_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _8989_ (.A1(_0849_),
    .A2(_0426_),
    .Z(_4029_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _8990_ (.I(_0854_),
    .Z(_4030_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _8991_ (.I0(_4029_),
    .I1(_0360_),
    .S(_4030_),
    .Z(_4031_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _8992_ (.A1(_2794_),
    .A2(_0342_),
    .A3(_4031_),
    .ZN(_4032_));
 gf180mcu_fd_sc_mcu7t5v0__or3_1 _8993_ (.A1(_4010_),
    .A2(_4028_),
    .A3(_4032_),
    .Z(_4033_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _8994_ (.A1(_1087_),
    .A2(_1287_),
    .ZN(_4034_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _8995_ (.A1(_1287_),
    .A2(_4033_),
    .B1(_4034_),
    .B2(_0526_),
    .C(_3199_),
    .ZN(_4035_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _8996_ (.A1(_3230_),
    .A2(_4029_),
    .ZN(_4036_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _8997_ (.A1(_4027_),
    .A2(_4036_),
    .ZN(_4037_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _8998_ (.A1(_2223_),
    .A2(_4027_),
    .B1(_4035_),
    .B2(_4037_),
    .ZN(_4038_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _8999_ (.A1(_3189_),
    .A2(_4038_),
    .ZN(_0272_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _9000_ (.A1(_3492_),
    .A2(_3122_),
    .B(_4026_),
    .ZN(_4039_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _9001_ (.A1(_4479_),
    .A2(_0624_),
    .ZN(_4040_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _9002_ (.I(_3122_),
    .ZN(_4041_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _9003_ (.A1(_1921_),
    .A2(_1640_),
    .ZN(_4042_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_1 _9004_ (.A1(_4042_),
    .A2(_4030_),
    .B1(_1009_),
    .B2(_3123_),
    .C(_0619_),
    .ZN(_4043_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _9005_ (.A1(_2635_),
    .A2(_3266_),
    .B(_4041_),
    .C(_4043_),
    .ZN(_4044_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _9006_ (.A1(_4040_),
    .A2(_4034_),
    .B1(_4044_),
    .B2(_1287_),
    .C(_3230_),
    .ZN(_4045_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _9007_ (.A1(_3230_),
    .A2(_4040_),
    .B(_4045_),
    .ZN(_4046_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _9008_ (.A1(_4463_),
    .A2(_4039_),
    .B(_1634_),
    .ZN(_4047_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _9009_ (.A1(_4039_),
    .A2(_4046_),
    .B(_4047_),
    .ZN(_0273_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_1 _9010_ (.A1(_3214_),
    .A2(_1551_),
    .A3(_3126_),
    .A4(_1249_),
    .ZN(_4048_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _9011_ (.A1(_4026_),
    .A2(_4048_),
    .ZN(_4049_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _9012_ (.A1(_0620_),
    .A2(_4030_),
    .ZN(_4050_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _9013_ (.A1(_4050_),
    .A2(_3113_),
    .B1(_3114_),
    .B2(_1296_),
    .ZN(_4051_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _9014_ (.A1(_0621_),
    .A2(_4030_),
    .A3(_3216_),
    .ZN(_4052_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _9015_ (.A1(_3136_),
    .A2(_3216_),
    .B(_1589_),
    .ZN(_4053_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _9016_ (.A1(_3492_),
    .A2(_4051_),
    .B1(_4052_),
    .B2(_4053_),
    .ZN(_4054_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _9017_ (.A1(_1589_),
    .A2(_4049_),
    .ZN(_4055_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _9018_ (.A1(_4049_),
    .A2(_4054_),
    .B(_4055_),
    .C(_3742_),
    .ZN(_0274_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _9019_ (.A1(_1517_),
    .A2(_1622_),
    .A3(_1624_),
    .ZN(_4056_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _9020_ (.A1(_0553_),
    .A2(_1364_),
    .ZN(_4057_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _9021_ (.A1(_4491_),
    .A2(_3268_),
    .A3(_2404_),
    .A4(_4057_),
    .ZN(_4058_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _9022_ (.A1(_2776_),
    .A2(_1317_),
    .B(_3282_),
    .C(_4058_),
    .ZN(_4059_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _9023_ (.A1(_1359_),
    .A2(_4059_),
    .ZN(_4060_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _9024_ (.A1(_1234_),
    .A2(_1233_),
    .A3(_1466_),
    .ZN(_4061_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _9025_ (.A1(_2395_),
    .A2(_1264_),
    .ZN(_4062_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _9026_ (.A1(_1463_),
    .A2(_4061_),
    .A3(_4062_),
    .ZN(_4063_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_2 _9027_ (.A1(_1475_),
    .A2(_2447_),
    .A3(_4060_),
    .A4(_4063_),
    .ZN(_4064_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _9028_ (.A1(_0855_),
    .A2(_4017_),
    .Z(_4065_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _9029_ (.A1(_4365_),
    .A2(_1251_),
    .ZN(_4066_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _9030_ (.A1(_3827_),
    .A2(_0516_),
    .B(_2631_),
    .C(_1034_),
    .ZN(_4067_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _9031_ (.A1(_2450_),
    .A2(_3074_),
    .A3(_4067_),
    .ZN(_4068_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _9032_ (.A1(_1163_),
    .A2(_4066_),
    .B(_4068_),
    .ZN(_4069_));
 gf180mcu_fd_sc_mcu7t5v0__and4_1 _9033_ (.A1(_1476_),
    .A2(_4064_),
    .A3(_4065_),
    .A4(_4069_),
    .Z(_4070_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _9034_ (.A1(_1291_),
    .A2(_4056_),
    .B(_4070_),
    .ZN(_4071_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _9035_ (.A1(_4430_),
    .A2(_1527_),
    .Z(_4072_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _9036_ (.A1(_4072_),
    .A2(_1290_),
    .B(_1520_),
    .ZN(_4073_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _9037_ (.A1(_1627_),
    .A2(_0566_),
    .B1(_3141_),
    .B2(_4073_),
    .ZN(_4074_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _9038_ (.A1(_3851_),
    .A2(_4074_),
    .B(_3868_),
    .ZN(_4075_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _9039_ (.A1(_3088_),
    .A2(_0570_),
    .ZN(_4076_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _9040_ (.A1(_1451_),
    .A2(_4075_),
    .B(_4071_),
    .C(_4076_),
    .ZN(_4077_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _9041_ (.A1(_1595_),
    .A2(_4071_),
    .B(_4077_),
    .C(_3742_),
    .ZN(_0275_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _9042_ (.A1(_1691_),
    .A2(_4056_),
    .B(_4070_),
    .ZN(_4078_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _9043_ (.A1(_0299_),
    .A2(_0320_),
    .Z(_4079_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _9044_ (.A1(_0299_),
    .A2(_0319_),
    .B(_4343_),
    .ZN(_4080_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _9045_ (.A1(_4335_),
    .A2(_4080_),
    .ZN(_4081_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _9046_ (.A1(_0421_),
    .A2(_0451_),
    .B1(_4079_),
    .B2(_4081_),
    .ZN(_4082_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _9047_ (.A1(_0421_),
    .A2(_0451_),
    .B1(_0467_),
    .B2(_0475_),
    .ZN(_4083_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _9048_ (.A1(_0561_),
    .A2(_0569_),
    .B1(_4082_),
    .B2(_4083_),
    .ZN(_4084_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _9049_ (.A1(_0467_),
    .A2(_0476_),
    .B(_4084_),
    .ZN(_4085_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _9050_ (.A1(_0561_),
    .A2(_0569_),
    .B1(_0653_),
    .B2(_0661_),
    .C(_4085_),
    .ZN(_4086_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _9051_ (.A1(_0653_),
    .A2(_0661_),
    .B1(_0732_),
    .B2(_0739_),
    .ZN(_4087_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _9052_ (.A1(_0732_),
    .A2(_0739_),
    .ZN(_4088_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_1 _9053_ (.A1(_0821_),
    .A2(_1431_),
    .B1(_4086_),
    .B2(_4087_),
    .C(_4088_),
    .ZN(_4089_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _9054_ (.A1(_0821_),
    .A2(_1431_),
    .B(_1518_),
    .ZN(_4090_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _9055_ (.A1(_4072_),
    .A2(_3113_),
    .B(_1519_),
    .ZN(_4091_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _9056_ (.A1(_1627_),
    .A2(_0818_),
    .B1(_3115_),
    .B2(_4091_),
    .C(_1628_),
    .ZN(_4092_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _9057_ (.A1(_3851_),
    .A2(_1100_),
    .B(_4092_),
    .ZN(_4093_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _9058_ (.A1(_4089_),
    .A2(_4090_),
    .B1(_4093_),
    .B2(_1576_),
    .C(_4078_),
    .ZN(_4094_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _9059_ (.A1(_4316_),
    .A2(_4078_),
    .B(_4094_),
    .C(_3742_),
    .ZN(_0276_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_1 _9060_ (.A1(_3106_),
    .A2(_1046_),
    .A3(_1244_),
    .A4(_2631_),
    .ZN(_4095_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _9061_ (.A1(_1575_),
    .A2(_4010_),
    .ZN(_4096_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _9062_ (.A1(_4064_),
    .A2(_4095_),
    .A3(_4096_),
    .ZN(_4097_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _9063_ (.A1(_1212_),
    .A2(_1431_),
    .Z(_4098_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _9064_ (.A1(_1518_),
    .A2(_0801_),
    .ZN(_4099_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _9065_ (.I(_4072_),
    .Z(_4100_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _9066_ (.A1(_4100_),
    .A2(_3128_),
    .B(_3127_),
    .ZN(_4101_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _9067_ (.A1(_4098_),
    .A2(_4099_),
    .B1(_4101_),
    .B2(_1576_),
    .C(_4097_),
    .ZN(_4102_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _9068_ (.A1(_3812_),
    .A2(_4097_),
    .B(_4102_),
    .C(_3249_),
    .ZN(_0277_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _9069_ (.A1(_2793_),
    .A2(_1469_),
    .ZN(_4103_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _9070_ (.A1(_3770_),
    .A2(_3268_),
    .A3(_4062_),
    .ZN(_4104_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_4 _9071_ (.A1(_1270_),
    .A2(_1274_),
    .A3(_4103_),
    .A4(_4104_),
    .ZN(_4105_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _9072_ (.A1(_2373_),
    .A2(_3144_),
    .B(_4105_),
    .ZN(_4106_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _9073_ (.A1(_1089_),
    .A2(_4106_),
    .ZN(_4107_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _9074_ (.I(_4105_),
    .Z(_4108_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _9075_ (.A1(_4100_),
    .A2(_3135_),
    .ZN(_4109_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _9076_ (.A1(_3138_),
    .A2(_4108_),
    .A3(_4109_),
    .ZN(_4110_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _9077_ (.A1(_4107_),
    .A2(_4110_),
    .B(_3619_),
    .ZN(_0278_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _9078_ (.A1(_3132_),
    .A2(_4105_),
    .ZN(_4111_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _9079_ (.A1(_4365_),
    .A2(_4111_),
    .ZN(_4112_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _9080_ (.I(_1622_),
    .Z(_4113_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _9081_ (.A1(_4113_),
    .A2(_4100_),
    .B(_3133_),
    .ZN(_4114_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _9082_ (.A1(_4108_),
    .A2(_4114_),
    .ZN(_4115_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _9083_ (.A1(_4112_),
    .A2(_4115_),
    .B(_3619_),
    .ZN(_0279_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _9084_ (.A1(_1552_),
    .A2(_3136_),
    .A3(_4100_),
    .ZN(_4116_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _9085_ (.A1(_1382_),
    .A2(_4113_),
    .B(_4116_),
    .ZN(_4117_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _9086_ (.A1(_4041_),
    .A2(_4108_),
    .B(\as2650.psl[1] ),
    .ZN(_4118_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _9087_ (.A1(_4108_),
    .A2(_4117_),
    .B(_4118_),
    .C(_3249_),
    .ZN(_0280_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _9088_ (.A1(_1523_),
    .A2(_0339_),
    .A3(_4062_),
    .ZN(_4119_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_1 _9089_ (.A1(_1319_),
    .A2(_2925_),
    .A3(_1245_),
    .A4(_4119_),
    .ZN(_4120_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _9090_ (.A1(_4065_),
    .A2(_4120_),
    .Z(_4121_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _9091_ (.I(_4121_),
    .Z(_4122_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _9092_ (.A1(_1706_),
    .A2(_4028_),
    .ZN(_4123_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _9093_ (.A1(_0944_),
    .A2(_4113_),
    .B(_4123_),
    .ZN(_4124_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _9094_ (.A1(_1588_),
    .A2(_4113_),
    .ZN(_4125_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _9095_ (.A1(_4125_),
    .A2(_4122_),
    .B(net27),
    .ZN(_4126_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _9096_ (.A1(_4122_),
    .A2(_4124_),
    .B(_4126_),
    .C(_3249_),
    .ZN(_0281_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _9097_ (.A1(_2373_),
    .A2(_3144_),
    .B(_4121_),
    .ZN(_4127_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _9098_ (.A1(\as2650.psu[4] ),
    .A2(_4127_),
    .ZN(_4128_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _9099_ (.A1(_1296_),
    .A2(_3137_),
    .B(_3135_),
    .ZN(_4129_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _9100_ (.A1(_4122_),
    .A2(_4129_),
    .ZN(_4130_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _9101_ (.A1(_4128_),
    .A2(_4130_),
    .B(_3619_),
    .ZN(_0282_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _9102_ (.A1(_3132_),
    .A2(_4121_),
    .ZN(_4131_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _9103_ (.A1(\as2650.psu[3] ),
    .A2(_4131_),
    .ZN(_4132_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _9104_ (.A1(_3133_),
    .A2(_4028_),
    .ZN(_4133_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _9105_ (.A1(_4122_),
    .A2(_4133_),
    .ZN(_4134_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _9106_ (.A1(_4132_),
    .A2(_4134_),
    .B(_1302_),
    .ZN(_0283_));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9107_ (.D(_0000_),
    .CLK(clknet_leaf_66_wb_clk_i),
    .Q(\as2650.r123[0][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9108_ (.D(_0001_),
    .CLK(clknet_leaf_68_wb_clk_i),
    .Q(\as2650.r123[0][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9109_ (.D(_0002_),
    .CLK(clknet_leaf_68_wb_clk_i),
    .Q(\as2650.r123[0][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9110_ (.D(_0003_),
    .CLK(clknet_leaf_68_wb_clk_i),
    .Q(\as2650.r123[0][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9111_ (.D(_0004_),
    .CLK(clknet_leaf_68_wb_clk_i),
    .Q(\as2650.r123[0][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9112_ (.D(_0005_),
    .CLK(clknet_leaf_68_wb_clk_i),
    .Q(\as2650.r123[0][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9113_ (.D(_0006_),
    .CLK(clknet_leaf_67_wb_clk_i),
    .Q(\as2650.r123[0][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9114_ (.D(_0007_),
    .CLK(clknet_leaf_67_wb_clk_i),
    .Q(\as2650.r123[0][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9115_ (.D(_0008_),
    .CLK(clknet_leaf_38_wb_clk_i),
    .Q(\as2650.stack[5][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9116_ (.D(_0009_),
    .CLK(clknet_leaf_42_wb_clk_i),
    .Q(\as2650.stack[5][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9117_ (.D(_0010_),
    .CLK(clknet_leaf_41_wb_clk_i),
    .Q(\as2650.stack[5][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9118_ (.D(_0011_),
    .CLK(clknet_leaf_39_wb_clk_i),
    .Q(\as2650.stack[5][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9119_ (.D(_0012_),
    .CLK(clknet_leaf_38_wb_clk_i),
    .Q(\as2650.stack[5][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9120_ (.D(_0013_),
    .CLK(clknet_leaf_38_wb_clk_i),
    .Q(\as2650.stack[5][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9121_ (.D(_0014_),
    .CLK(clknet_leaf_39_wb_clk_i),
    .Q(\as2650.stack[5][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9122_ (.D(_0015_),
    .CLK(clknet_leaf_42_wb_clk_i),
    .Q(\as2650.stack[5][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9123_ (.D(_0016_),
    .CLK(clknet_leaf_58_wb_clk_i),
    .Q(\as2650.stack[6][8] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9124_ (.D(_0017_),
    .CLK(clknet_leaf_57_wb_clk_i),
    .Q(\as2650.stack[6][9] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9125_ (.D(_0018_),
    .CLK(clknet_leaf_57_wb_clk_i),
    .Q(\as2650.stack[6][10] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9126_ (.D(_0019_),
    .CLK(clknet_leaf_59_wb_clk_i),
    .Q(\as2650.stack[6][11] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9127_ (.D(_0020_),
    .CLK(clknet_leaf_58_wb_clk_i),
    .Q(\as2650.stack[6][12] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9128_ (.D(_0021_),
    .CLK(clknet_leaf_58_wb_clk_i),
    .Q(\as2650.stack[6][13] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9129_ (.D(_0022_),
    .CLK(clknet_leaf_58_wb_clk_i),
    .Q(\as2650.stack[6][14] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9130_ (.D(_0023_),
    .CLK(clknet_leaf_58_wb_clk_i),
    .Q(\as2650.stack[5][8] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9131_ (.D(_0024_),
    .CLK(clknet_leaf_49_wb_clk_i),
    .Q(\as2650.stack[5][9] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9132_ (.D(_0025_),
    .CLK(clknet_leaf_56_wb_clk_i),
    .Q(\as2650.stack[5][10] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9133_ (.D(_0026_),
    .CLK(clknet_leaf_53_wb_clk_i),
    .Q(\as2650.stack[5][11] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9134_ (.D(_0027_),
    .CLK(clknet_leaf_56_wb_clk_i),
    .Q(\as2650.stack[5][12] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9135_ (.D(_0028_),
    .CLK(clknet_leaf_58_wb_clk_i),
    .Q(\as2650.stack[5][13] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9136_ (.D(_0029_),
    .CLK(clknet_leaf_58_wb_clk_i),
    .Q(\as2650.stack[5][14] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9137_ (.D(_0030_),
    .CLK(clknet_leaf_46_wb_clk_i),
    .Q(\as2650.r123_2[0][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9138_ (.D(_0031_),
    .CLK(clknet_leaf_46_wb_clk_i),
    .Q(\as2650.r123_2[0][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9139_ (.D(_0032_),
    .CLK(clknet_leaf_46_wb_clk_i),
    .Q(\as2650.r123_2[0][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9140_ (.D(_0033_),
    .CLK(clknet_leaf_46_wb_clk_i),
    .Q(\as2650.r123_2[0][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9141_ (.D(_0034_),
    .CLK(clknet_leaf_67_wb_clk_i),
    .Q(\as2650.r123_2[0][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9142_ (.D(_0035_),
    .CLK(clknet_leaf_67_wb_clk_i),
    .Q(\as2650.r123_2[0][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9143_ (.D(_0036_),
    .CLK(clknet_leaf_67_wb_clk_i),
    .Q(\as2650.r123_2[0][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9144_ (.D(_0037_),
    .CLK(clknet_leaf_66_wb_clk_i),
    .Q(\as2650.r123_2[0][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9145_ (.D(_0038_),
    .CLK(clknet_leaf_6_wb_clk_i),
    .Q(\as2650.psu[5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9146_ (.D(_0039_),
    .CLK(clknet_leaf_15_wb_clk_i),
    .Q(net41));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9147_ (.D(_0040_),
    .CLK(clknet_leaf_15_wb_clk_i),
    .Q(net42));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9148_ (.D(_0041_),
    .CLK(clknet_leaf_15_wb_clk_i),
    .Q(net43));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9149_ (.D(_0042_),
    .CLK(clknet_leaf_15_wb_clk_i),
    .Q(net44));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9150_ (.D(_0043_),
    .CLK(clknet_leaf_15_wb_clk_i),
    .Q(net45));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9151_ (.D(_0044_),
    .CLK(clknet_leaf_15_wb_clk_i),
    .Q(net19));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9152_ (.D(_0045_),
    .CLK(clknet_leaf_16_wb_clk_i),
    .Q(net20));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9153_ (.D(_0046_),
    .CLK(clknet_leaf_16_wb_clk_i),
    .Q(net21));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9154_ (.D(_0047_),
    .CLK(clknet_leaf_57_wb_clk_i),
    .Q(\as2650.stack[4][8] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9155_ (.D(_0048_),
    .CLK(clknet_leaf_57_wb_clk_i),
    .Q(\as2650.stack[4][9] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9156_ (.D(_0049_),
    .CLK(clknet_leaf_56_wb_clk_i),
    .Q(\as2650.stack[4][10] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9157_ (.D(_0050_),
    .CLK(clknet_leaf_57_wb_clk_i),
    .Q(\as2650.stack[4][11] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9158_ (.D(_0051_),
    .CLK(clknet_leaf_56_wb_clk_i),
    .Q(\as2650.stack[4][12] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9159_ (.D(_0052_),
    .CLK(clknet_leaf_58_wb_clk_i),
    .Q(\as2650.stack[4][13] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9160_ (.D(_0053_),
    .CLK(clknet_leaf_58_wb_clk_i),
    .Q(\as2650.stack[4][14] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9161_ (.D(_0054_),
    .CLK(clknet_3_4_0_wb_clk_i),
    .Q(\as2650.psl[6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9162_ (.D(_0055_),
    .CLK(clknet_leaf_45_wb_clk_i),
    .Q(\as2650.psl[7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9163_ (.D(_0056_),
    .CLK(clknet_leaf_48_wb_clk_i),
    .Q(\as2650.stack[3][8] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9164_ (.D(_0057_),
    .CLK(clknet_leaf_48_wb_clk_i),
    .Q(\as2650.stack[3][9] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9165_ (.D(_0058_),
    .CLK(clknet_leaf_48_wb_clk_i),
    .Q(\as2650.stack[3][10] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9166_ (.D(_0059_),
    .CLK(clknet_leaf_48_wb_clk_i),
    .Q(\as2650.stack[3][11] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9167_ (.D(_0060_),
    .CLK(clknet_leaf_49_wb_clk_i),
    .Q(\as2650.stack[3][12] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9168_ (.D(_0061_),
    .CLK(clknet_leaf_48_wb_clk_i),
    .Q(\as2650.stack[3][13] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9169_ (.D(_0062_),
    .CLK(clknet_leaf_48_wb_clk_i),
    .Q(\as2650.stack[3][14] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9170_ (.D(_0063_),
    .CLK(clknet_leaf_60_wb_clk_i),
    .Q(\as2650.stack[2][8] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9171_ (.D(_0064_),
    .CLK(clknet_leaf_60_wb_clk_i),
    .Q(\as2650.stack[2][9] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9172_ (.D(_0065_),
    .CLK(clknet_leaf_60_wb_clk_i),
    .Q(\as2650.stack[2][10] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9173_ (.D(_0066_),
    .CLK(clknet_leaf_60_wb_clk_i),
    .Q(\as2650.stack[2][11] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9174_ (.D(_0067_),
    .CLK(clknet_leaf_60_wb_clk_i),
    .Q(\as2650.stack[2][12] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9175_ (.D(_0068_),
    .CLK(clknet_leaf_60_wb_clk_i),
    .Q(\as2650.stack[2][13] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9176_ (.D(_0069_),
    .CLK(clknet_leaf_59_wb_clk_i),
    .Q(\as2650.stack[2][14] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9177_ (.D(_0070_),
    .CLK(clknet_leaf_71_wb_clk_i),
    .Q(\as2650.ins_reg[0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9178_ (.D(_0071_),
    .CLK(clknet_leaf_73_wb_clk_i),
    .Q(\as2650.ins_reg[1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9179_ (.D(_0072_),
    .CLK(clknet_leaf_9_wb_clk_i),
    .Q(\as2650.ins_reg[2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9180_ (.D(_0073_),
    .CLK(clknet_leaf_6_wb_clk_i),
    .Q(\as2650.ins_reg[5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9181_ (.D(_0074_),
    .CLK(clknet_leaf_8_wb_clk_i),
    .Q(\as2650.ins_reg[6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9182_ (.D(_0075_),
    .CLK(clknet_leaf_8_wb_clk_i),
    .Q(\as2650.ins_reg[7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9183_ (.D(_0076_),
    .CLK(clknet_leaf_74_wb_clk_i),
    .Q(\as2650.r123_2[1][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9184_ (.D(_0077_),
    .CLK(clknet_leaf_69_wb_clk_i),
    .Q(\as2650.r123_2[1][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9185_ (.D(_0078_),
    .CLK(clknet_leaf_73_wb_clk_i),
    .Q(\as2650.r123_2[1][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9186_ (.D(_0079_),
    .CLK(clknet_leaf_73_wb_clk_i),
    .Q(\as2650.r123_2[1][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9187_ (.D(_0080_),
    .CLK(clknet_leaf_65_wb_clk_i),
    .Q(\as2650.r123_2[1][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9188_ (.D(_0081_),
    .CLK(clknet_leaf_69_wb_clk_i),
    .Q(\as2650.r123_2[1][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9189_ (.D(_0082_),
    .CLK(clknet_leaf_65_wb_clk_i),
    .Q(\as2650.r123_2[1][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9190_ (.D(_0083_),
    .CLK(clknet_leaf_65_wb_clk_i),
    .Q(\as2650.r123_2[1][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9191_ (.D(_0084_),
    .CLK(clknet_leaf_47_wb_clk_i),
    .Q(\as2650.stack[1][8] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9192_ (.D(_0085_),
    .CLK(clknet_leaf_48_wb_clk_i),
    .Q(\as2650.stack[1][9] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9193_ (.D(_0086_),
    .CLK(clknet_leaf_48_wb_clk_i),
    .Q(\as2650.stack[1][10] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9194_ (.D(_0087_),
    .CLK(clknet_leaf_48_wb_clk_i),
    .Q(\as2650.stack[1][11] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9195_ (.D(_0088_),
    .CLK(clknet_leaf_47_wb_clk_i),
    .Q(\as2650.stack[1][12] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9196_ (.D(_0089_),
    .CLK(clknet_leaf_47_wb_clk_i),
    .Q(\as2650.stack[1][13] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9197_ (.D(_0090_),
    .CLK(clknet_leaf_47_wb_clk_i),
    .Q(\as2650.stack[1][14] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9198_ (.D(_0091_),
    .CLK(clknet_leaf_46_wb_clk_i),
    .Q(\as2650.stack[0][8] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9199_ (.D(_0092_),
    .CLK(clknet_leaf_47_wb_clk_i),
    .Q(\as2650.stack[0][9] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9200_ (.D(_0093_),
    .CLK(clknet_leaf_60_wb_clk_i),
    .Q(\as2650.stack[0][10] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9201_ (.D(_0094_),
    .CLK(clknet_leaf_60_wb_clk_i),
    .Q(\as2650.stack[0][11] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9202_ (.D(_0095_),
    .CLK(clknet_leaf_47_wb_clk_i),
    .Q(\as2650.stack[0][12] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9203_ (.D(_0096_),
    .CLK(clknet_leaf_47_wb_clk_i),
    .Q(\as2650.stack[0][13] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9204_ (.D(_0097_),
    .CLK(clknet_leaf_46_wb_clk_i),
    .Q(\as2650.stack[0][14] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9205_ (.D(_0098_),
    .CLK(clknet_leaf_74_wb_clk_i),
    .Q(\as2650.r123_2[2][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9206_ (.D(_0099_),
    .CLK(clknet_leaf_73_wb_clk_i),
    .Q(\as2650.r123_2[2][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9207_ (.D(_0100_),
    .CLK(clknet_leaf_77_wb_clk_i),
    .Q(\as2650.r123_2[2][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9208_ (.D(_0101_),
    .CLK(clknet_leaf_77_wb_clk_i),
    .Q(\as2650.r123_2[2][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9209_ (.D(_0102_),
    .CLK(clknet_leaf_75_wb_clk_i),
    .Q(\as2650.r123_2[2][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9210_ (.D(_0103_),
    .CLK(clknet_leaf_77_wb_clk_i),
    .Q(\as2650.r123_2[2][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9211_ (.D(_0104_),
    .CLK(clknet_leaf_76_wb_clk_i),
    .Q(\as2650.r123_2[2][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9212_ (.D(_0105_),
    .CLK(clknet_leaf_75_wb_clk_i),
    .Q(\as2650.r123_2[2][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9213_ (.D(_0106_),
    .CLK(clknet_leaf_56_wb_clk_i),
    .Q(\as2650.stack[2][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9214_ (.D(_0107_),
    .CLK(clknet_leaf_41_wb_clk_i),
    .Q(\as2650.stack[2][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9215_ (.D(_0108_),
    .CLK(clknet_leaf_41_wb_clk_i),
    .Q(\as2650.stack[2][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9216_ (.D(_0109_),
    .CLK(clknet_leaf_41_wb_clk_i),
    .Q(\as2650.stack[2][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9217_ (.D(_0110_),
    .CLK(clknet_leaf_53_wb_clk_i),
    .Q(\as2650.stack[2][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9218_ (.D(_0111_),
    .CLK(clknet_leaf_56_wb_clk_i),
    .Q(\as2650.stack[2][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9219_ (.D(_0112_),
    .CLK(clknet_leaf_54_wb_clk_i),
    .Q(\as2650.stack[2][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9220_ (.D(_0113_),
    .CLK(clknet_leaf_40_wb_clk_i),
    .Q(\as2650.stack[2][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9221_ (.D(_0114_),
    .CLK(clknet_leaf_37_wb_clk_i),
    .Q(\as2650.stack[4][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9222_ (.D(_0115_),
    .CLK(clknet_leaf_40_wb_clk_i),
    .Q(\as2650.stack[4][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9223_ (.D(_0116_),
    .CLK(clknet_leaf_40_wb_clk_i),
    .Q(\as2650.stack[4][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9224_ (.D(_0117_),
    .CLK(clknet_leaf_39_wb_clk_i),
    .Q(\as2650.stack[4][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9225_ (.D(_0118_),
    .CLK(clknet_leaf_55_wb_clk_i),
    .Q(\as2650.stack[4][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9226_ (.D(_0119_),
    .CLK(clknet_leaf_37_wb_clk_i),
    .Q(\as2650.stack[4][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9227_ (.D(_0120_),
    .CLK(clknet_leaf_36_wb_clk_i),
    .Q(\as2650.stack[4][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9228_ (.D(_0121_),
    .CLK(clknet_leaf_40_wb_clk_i),
    .Q(\as2650.stack[4][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9229_ (.D(_0122_),
    .CLK(clknet_leaf_62_wb_clk_i),
    .Q(\as2650.r123_2[3][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9230_ (.D(_0123_),
    .CLK(clknet_leaf_61_wb_clk_i),
    .Q(\as2650.r123_2[3][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9231_ (.D(_0124_),
    .CLK(clknet_leaf_61_wb_clk_i),
    .Q(\as2650.r123_2[3][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9232_ (.D(_0125_),
    .CLK(clknet_leaf_63_wb_clk_i),
    .Q(\as2650.r123_2[3][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9233_ (.D(_0126_),
    .CLK(clknet_3_0_0_wb_clk_i),
    .Q(\as2650.r123_2[3][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9234_ (.D(_0127_),
    .CLK(clknet_leaf_62_wb_clk_i),
    .Q(\as2650.r123_2[3][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9235_ (.D(_0128_),
    .CLK(clknet_leaf_62_wb_clk_i),
    .Q(\as2650.r123_2[3][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9236_ (.D(_0129_),
    .CLK(clknet_leaf_64_wb_clk_i),
    .Q(\as2650.r123_2[3][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9237_ (.D(_0130_),
    .CLK(clknet_leaf_55_wb_clk_i),
    .Q(\as2650.stack[1][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9238_ (.D(_0131_),
    .CLK(clknet_leaf_39_wb_clk_i),
    .Q(\as2650.stack[1][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9239_ (.D(_0132_),
    .CLK(clknet_leaf_39_wb_clk_i),
    .Q(\as2650.stack[1][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9240_ (.D(_0133_),
    .CLK(clknet_leaf_38_wb_clk_i),
    .Q(\as2650.stack[1][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9241_ (.D(_0134_),
    .CLK(clknet_leaf_55_wb_clk_i),
    .Q(\as2650.stack[1][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9242_ (.D(_0135_),
    .CLK(clknet_leaf_55_wb_clk_i),
    .Q(\as2650.stack[1][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9243_ (.D(_0136_),
    .CLK(clknet_leaf_55_wb_clk_i),
    .Q(\as2650.stack[1][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9244_ (.D(_0137_),
    .CLK(clknet_leaf_39_wb_clk_i),
    .Q(\as2650.stack[1][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9245_ (.D(_0138_),
    .CLK(clknet_3_0_0_wb_clk_i),
    .Q(\as2650.r123[3][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9246_ (.D(_0139_),
    .CLK(clknet_leaf_62_wb_clk_i),
    .Q(\as2650.r123[3][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9247_ (.D(_0140_),
    .CLK(clknet_leaf_62_wb_clk_i),
    .Q(\as2650.r123[3][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9248_ (.D(_0141_),
    .CLK(clknet_leaf_63_wb_clk_i),
    .Q(\as2650.r123[3][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9249_ (.D(_0142_),
    .CLK(clknet_3_1_0_wb_clk_i),
    .Q(\as2650.r123[3][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9250_ (.D(_0143_),
    .CLK(clknet_leaf_64_wb_clk_i),
    .Q(\as2650.r123[3][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9251_ (.D(_0144_),
    .CLK(clknet_leaf_63_wb_clk_i),
    .Q(\as2650.r123[3][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9252_ (.D(_0145_),
    .CLK(clknet_leaf_63_wb_clk_i),
    .Q(\as2650.r123[3][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9253_ (.D(_0146_),
    .CLK(clknet_leaf_55_wb_clk_i),
    .Q(\as2650.stack[3][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9254_ (.D(_0147_),
    .CLK(clknet_leaf_50_wb_clk_i),
    .Q(\as2650.stack[3][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9255_ (.D(_0148_),
    .CLK(clknet_leaf_50_wb_clk_i),
    .Q(\as2650.stack[3][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9256_ (.D(_0149_),
    .CLK(clknet_leaf_44_wb_clk_i),
    .Q(\as2650.stack[3][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9257_ (.D(_0150_),
    .CLK(clknet_leaf_55_wb_clk_i),
    .Q(\as2650.stack[3][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9258_ (.D(_0151_),
    .CLK(clknet_leaf_56_wb_clk_i),
    .Q(\as2650.stack[3][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9259_ (.D(_0152_),
    .CLK(clknet_leaf_55_wb_clk_i),
    .Q(\as2650.stack[3][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9260_ (.D(_0153_),
    .CLK(clknet_leaf_50_wb_clk_i),
    .Q(\as2650.stack[3][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9261_ (.D(_0154_),
    .CLK(clknet_leaf_54_wb_clk_i),
    .Q(\as2650.stack[0][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9262_ (.D(_0155_),
    .CLK(clknet_leaf_51_wb_clk_i),
    .Q(\as2650.stack[0][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9263_ (.D(_0156_),
    .CLK(clknet_leaf_52_wb_clk_i),
    .Q(\as2650.stack[0][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9264_ (.D(_0157_),
    .CLK(clknet_leaf_52_wb_clk_i),
    .Q(\as2650.stack[0][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9265_ (.D(_0158_),
    .CLK(clknet_leaf_54_wb_clk_i),
    .Q(\as2650.stack[0][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9266_ (.D(_0159_),
    .CLK(clknet_leaf_54_wb_clk_i),
    .Q(\as2650.stack[0][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9267_ (.D(_0160_),
    .CLK(clknet_leaf_54_wb_clk_i),
    .Q(\as2650.stack[0][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9268_ (.D(_0161_),
    .CLK(clknet_leaf_52_wb_clk_i),
    .Q(\as2650.stack[0][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9269_ (.D(_0162_),
    .CLK(clknet_leaf_14_wb_clk_i),
    .Q(\as2650.addr_buff[0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9270_ (.D(_0163_),
    .CLK(clknet_leaf_12_wb_clk_i),
    .Q(\as2650.addr_buff[1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9271_ (.D(_0164_),
    .CLK(clknet_leaf_14_wb_clk_i),
    .Q(\as2650.addr_buff[2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9272_ (.D(_0165_),
    .CLK(clknet_leaf_12_wb_clk_i),
    .Q(\as2650.addr_buff[3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9273_ (.D(_0166_),
    .CLK(clknet_leaf_12_wb_clk_i),
    .Q(\as2650.addr_buff[4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9274_ (.D(_0167_),
    .CLK(clknet_leaf_11_wb_clk_i),
    .Q(\as2650.addr_buff[5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9275_ (.D(_0168_),
    .CLK(clknet_leaf_11_wb_clk_i),
    .Q(\as2650.addr_buff[6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9276_ (.D(_0169_),
    .CLK(clknet_3_2_0_wb_clk_i),
    .Q(\as2650.addr_buff[7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9277_ (.D(_0170_),
    .CLK(clknet_leaf_20_wb_clk_i),
    .Q(net24));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9278_ (.D(_0171_),
    .CLK(clknet_leaf_20_wb_clk_i),
    .Q(net22));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9279_ (.D(_0172_),
    .CLK(clknet_3_3_0_wb_clk_i),
    .Q(net23));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9280_ (.D(_0173_),
    .CLK(clknet_leaf_26_wb_clk_i),
    .Q(net28));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9281_ (.D(_0174_),
    .CLK(clknet_leaf_26_wb_clk_i),
    .Q(net29));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9282_ (.D(_0175_),
    .CLK(clknet_leaf_26_wb_clk_i),
    .Q(net30));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9283_ (.D(_0176_),
    .CLK(clknet_leaf_26_wb_clk_i),
    .Q(net31));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9284_ (.D(_0177_),
    .CLK(clknet_leaf_26_wb_clk_i),
    .Q(net32));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9285_ (.D(_0178_),
    .CLK(clknet_leaf_27_wb_clk_i),
    .Q(net33));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9286_ (.D(_0179_),
    .CLK(clknet_leaf_27_wb_clk_i),
    .Q(net34));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9287_ (.D(_0180_),
    .CLK(clknet_leaf_27_wb_clk_i),
    .Q(net35));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9288_ (.D(_0181_),
    .CLK(clknet_leaf_27_wb_clk_i),
    .Q(net36));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9289_ (.D(_0182_),
    .CLK(clknet_leaf_28_wb_clk_i),
    .Q(net37));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9290_ (.D(_0183_),
    .CLK(clknet_leaf_28_wb_clk_i),
    .Q(net38));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9291_ (.D(_0184_),
    .CLK(clknet_leaf_31_wb_clk_i),
    .Q(net39));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9292_ (.D(_0185_),
    .CLK(clknet_leaf_31_wb_clk_i),
    .Q(net40));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9293_ (.D(_0186_),
    .CLK(clknet_leaf_20_wb_clk_i),
    .Q(net26));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9294_ (.D(_0187_),
    .CLK(clknet_leaf_25_wb_clk_i),
    .Q(net25));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9295_ (.D(_0188_),
    .CLK(clknet_leaf_11_wb_clk_i),
    .Q(\as2650.idx_ctrl[0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9296_ (.D(_0189_),
    .CLK(clknet_leaf_11_wb_clk_i),
    .Q(\as2650.idx_ctrl[1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9297_ (.D(_0190_),
    .CLK(clknet_leaf_3_wb_clk_i),
    .Q(\as2650.holding_reg[0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9298_ (.D(_0191_),
    .CLK(clknet_leaf_2_wb_clk_i),
    .Q(\as2650.holding_reg[1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9299_ (.D(_0192_),
    .CLK(clknet_leaf_1_wb_clk_i),
    .Q(\as2650.holding_reg[2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9300_ (.D(_0193_),
    .CLK(clknet_leaf_1_wb_clk_i),
    .Q(\as2650.holding_reg[3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9301_ (.D(_0194_),
    .CLK(clknet_leaf_1_wb_clk_i),
    .Q(\as2650.holding_reg[4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9302_ (.D(_0195_),
    .CLK(clknet_leaf_1_wb_clk_i),
    .Q(\as2650.holding_reg[5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9303_ (.D(_0196_),
    .CLK(clknet_leaf_2_wb_clk_i),
    .Q(\as2650.holding_reg[6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9304_ (.D(_0197_),
    .CLK(clknet_3_0_0_wb_clk_i),
    .Q(\as2650.holding_reg[7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9305_ (.D(_0198_),
    .CLK(clknet_3_3_0_wb_clk_i),
    .Q(\as2650.halted ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9306_ (.D(_0199_),
    .CLK(clknet_leaf_23_wb_clk_i),
    .Q(\as2650.cycle[0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9307_ (.D(_0200_),
    .CLK(clknet_leaf_23_wb_clk_i),
    .Q(\as2650.cycle[1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9308_ (.D(_0201_),
    .CLK(clknet_leaf_18_wb_clk_i),
    .Q(\as2650.cycle[2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_2 _9309_ (.D(_0202_),
    .CLK(clknet_leaf_16_wb_clk_i),
    .Q(\as2650.cycle[3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9310_ (.D(_0203_),
    .CLK(clknet_leaf_18_wb_clk_i),
    .Q(\as2650.cycle[4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_2 _9311_ (.D(_0204_),
    .CLK(clknet_3_3_0_wb_clk_i),
    .Q(\as2650.cycle[5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9312_ (.D(_0205_),
    .CLK(clknet_leaf_18_wb_clk_i),
    .Q(\as2650.cycle[6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9313_ (.D(_0206_),
    .CLK(clknet_leaf_18_wb_clk_i),
    .Q(\as2650.cycle[7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9314_ (.D(_0207_),
    .CLK(clknet_leaf_9_wb_clk_i),
    .Q(\as2650.psu[7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9315_ (.D(_0208_),
    .CLK(clknet_leaf_24_wb_clk_i),
    .Q(\as2650.pc[0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9316_ (.D(_0209_),
    .CLK(clknet_3_2_0_wb_clk_i),
    .Q(\as2650.pc[1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9317_ (.D(_0210_),
    .CLK(clknet_leaf_25_wb_clk_i),
    .Q(\as2650.pc[2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9318_ (.D(_0211_),
    .CLK(clknet_leaf_30_wb_clk_i),
    .Q(\as2650.pc[3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9319_ (.D(_0212_),
    .CLK(clknet_3_6_0_wb_clk_i),
    .Q(\as2650.pc[4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9320_ (.D(_0213_),
    .CLK(clknet_leaf_31_wb_clk_i),
    .Q(\as2650.pc[5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9321_ (.D(_0214_),
    .CLK(clknet_leaf_31_wb_clk_i),
    .Q(\as2650.pc[6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9322_ (.D(_0215_),
    .CLK(clknet_leaf_29_wb_clk_i),
    .Q(\as2650.pc[7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9323_ (.D(_0216_),
    .CLK(clknet_leaf_24_wb_clk_i),
    .Q(\as2650.pc[8] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9324_ (.D(_0217_),
    .CLK(clknet_leaf_29_wb_clk_i),
    .Q(\as2650.pc[9] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9325_ (.D(_0218_),
    .CLK(clknet_leaf_30_wb_clk_i),
    .Q(\as2650.pc[10] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9326_ (.D(_0219_),
    .CLK(clknet_3_6_0_wb_clk_i),
    .Q(\as2650.pc[11] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9327_ (.D(_0220_),
    .CLK(clknet_3_7_0_wb_clk_i),
    .Q(\as2650.pc[12] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9328_ (.D(_0221_),
    .CLK(clknet_3_7_0_wb_clk_i),
    .Q(\as2650.pc[13] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9329_ (.D(_0222_),
    .CLK(clknet_3_6_0_wb_clk_i),
    .Q(\as2650.pc[14] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9330_ (.D(_0223_),
    .CLK(clknet_leaf_80_wb_clk_i),
    .Q(\as2650.r0[0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9331_ (.D(_0224_),
    .CLK(clknet_leaf_80_wb_clk_i),
    .Q(\as2650.r0[1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9332_ (.D(_0225_),
    .CLK(clknet_leaf_80_wb_clk_i),
    .Q(\as2650.r0[2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9333_ (.D(_0226_),
    .CLK(clknet_leaf_80_wb_clk_i),
    .Q(\as2650.r0[3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9334_ (.D(_0227_),
    .CLK(clknet_leaf_80_wb_clk_i),
    .Q(\as2650.r0[4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9335_ (.D(_0228_),
    .CLK(clknet_leaf_80_wb_clk_i),
    .Q(\as2650.r0[5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9336_ (.D(_0229_),
    .CLK(clknet_3_0_0_wb_clk_i),
    .Q(\as2650.r0[6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9337_ (.D(_0230_),
    .CLK(clknet_leaf_77_wb_clk_i),
    .Q(\as2650.r0[7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9338_ (.D(_0231_),
    .CLK(clknet_leaf_39_wb_clk_i),
    .Q(\as2650.stack[6][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9339_ (.D(_0232_),
    .CLK(clknet_leaf_51_wb_clk_i),
    .Q(\as2650.stack[6][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9340_ (.D(_0233_),
    .CLK(clknet_leaf_50_wb_clk_i),
    .Q(\as2650.stack[6][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9341_ (.D(_0234_),
    .CLK(clknet_leaf_51_wb_clk_i),
    .Q(\as2650.stack[6][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9342_ (.D(_0235_),
    .CLK(clknet_leaf_38_wb_clk_i),
    .Q(\as2650.stack[6][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9343_ (.D(_0236_),
    .CLK(clknet_leaf_38_wb_clk_i),
    .Q(\as2650.stack[6][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9344_ (.D(_0237_),
    .CLK(clknet_leaf_37_wb_clk_i),
    .Q(\as2650.stack[6][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9345_ (.D(_0238_),
    .CLK(clknet_leaf_52_wb_clk_i),
    .Q(\as2650.stack[6][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9346_ (.D(_0239_),
    .CLK(clknet_leaf_37_wb_clk_i),
    .Q(\as2650.stack[7][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9347_ (.D(_0240_),
    .CLK(clknet_leaf_40_wb_clk_i),
    .Q(\as2650.stack[7][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9348_ (.D(_0241_),
    .CLK(clknet_leaf_41_wb_clk_i),
    .Q(\as2650.stack[7][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9349_ (.D(_0242_),
    .CLK(clknet_leaf_51_wb_clk_i),
    .Q(\as2650.stack[7][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9350_ (.D(_0243_),
    .CLK(clknet_leaf_36_wb_clk_i),
    .Q(\as2650.stack[7][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9351_ (.D(_0244_),
    .CLK(clknet_leaf_38_wb_clk_i),
    .Q(\as2650.stack[7][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9352_ (.D(_0245_),
    .CLK(clknet_leaf_38_wb_clk_i),
    .Q(\as2650.stack[7][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9353_ (.D(_0246_),
    .CLK(clknet_leaf_44_wb_clk_i),
    .Q(\as2650.stack[7][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9354_ (.D(_0247_),
    .CLK(clknet_leaf_59_wb_clk_i),
    .Q(\as2650.stack[7][8] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9355_ (.D(_0248_),
    .CLK(clknet_leaf_60_wb_clk_i),
    .Q(\as2650.stack[7][9] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9356_ (.D(_0249_),
    .CLK(clknet_leaf_59_wb_clk_i),
    .Q(\as2650.stack[7][10] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9357_ (.D(_0250_),
    .CLK(clknet_leaf_60_wb_clk_i),
    .Q(\as2650.stack[7][11] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9358_ (.D(_0251_),
    .CLK(clknet_leaf_59_wb_clk_i),
    .Q(\as2650.stack[7][12] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9359_ (.D(_0252_),
    .CLK(clknet_leaf_59_wb_clk_i),
    .Q(\as2650.stack[7][13] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9360_ (.D(_0253_),
    .CLK(clknet_leaf_59_wb_clk_i),
    .Q(\as2650.stack[7][14] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9361_ (.D(_0254_),
    .CLK(clknet_leaf_74_wb_clk_i),
    .Q(\as2650.r123[1][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9362_ (.D(_0255_),
    .CLK(clknet_leaf_69_wb_clk_i),
    .Q(\as2650.r123[1][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9363_ (.D(_0256_),
    .CLK(clknet_leaf_69_wb_clk_i),
    .Q(\as2650.r123[1][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9364_ (.D(_0257_),
    .CLK(clknet_leaf_73_wb_clk_i),
    .Q(\as2650.r123[1][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9365_ (.D(_0258_),
    .CLK(clknet_3_4_0_wb_clk_i),
    .Q(\as2650.r123[1][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9366_ (.D(_0259_),
    .CLK(clknet_leaf_68_wb_clk_i),
    .Q(\as2650.r123[1][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9367_ (.D(_0260_),
    .CLK(clknet_leaf_68_wb_clk_i),
    .Q(\as2650.r123[1][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9368_ (.D(_0261_),
    .CLK(clknet_leaf_65_wb_clk_i),
    .Q(\as2650.r123[1][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9369_ (.D(_0262_),
    .CLK(clknet_leaf_74_wb_clk_i),
    .Q(\as2650.r123[2][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9370_ (.D(_0263_),
    .CLK(clknet_leaf_76_wb_clk_i),
    .Q(\as2650.r123[2][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9371_ (.D(_0264_),
    .CLK(clknet_leaf_76_wb_clk_i),
    .Q(\as2650.r123[2][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9372_ (.D(_0265_),
    .CLK(clknet_leaf_76_wb_clk_i),
    .Q(\as2650.r123[2][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9373_ (.D(_0266_),
    .CLK(clknet_leaf_74_wb_clk_i),
    .Q(\as2650.r123[2][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9374_ (.D(_0267_),
    .CLK(clknet_leaf_77_wb_clk_i),
    .Q(\as2650.r123[2][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9375_ (.D(_0268_),
    .CLK(clknet_leaf_75_wb_clk_i),
    .Q(\as2650.r123[2][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9376_ (.D(_0269_),
    .CLK(clknet_leaf_74_wb_clk_i),
    .Q(\as2650.r123[2][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9377_ (.D(_0270_),
    .CLK(clknet_leaf_9_wb_clk_i),
    .Q(\as2650.ins_reg[3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9378_ (.D(_0271_),
    .CLK(clknet_leaf_8_wb_clk_i),
    .Q(\as2650.ins_reg[4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9379_ (.D(_0272_),
    .CLK(clknet_leaf_45_wb_clk_i),
    .Q(\as2650.psu[2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9380_ (.D(_0273_),
    .CLK(clknet_leaf_44_wb_clk_i),
    .Q(\as2650.psu[1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9381_ (.D(_0274_),
    .CLK(clknet_leaf_44_wb_clk_i),
    .Q(\as2650.psu[0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9382_ (.D(_0275_),
    .CLK(clknet_3_2_0_wb_clk_i),
    .Q(\as2650.psl[5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9383_ (.D(_0276_),
    .CLK(clknet_leaf_3_wb_clk_i),
    .Q(\as2650.carry ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9384_ (.D(_0277_),
    .CLK(clknet_leaf_3_wb_clk_i),
    .Q(\as2650.overflow ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9385_ (.D(_0278_),
    .CLK(clknet_leaf_71_wb_clk_i),
    .Q(\as2650.psl[4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9386_ (.D(_0279_),
    .CLK(clknet_leaf_3_wb_clk_i),
    .Q(\as2650.psl[3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9387_ (.D(_0280_),
    .CLK(clknet_leaf_5_wb_clk_i),
    .Q(\as2650.psl[1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9388_ (.D(_0281_),
    .CLK(clknet_3_1_0_wb_clk_i),
    .Q(net27));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9389_ (.D(_0282_),
    .CLK(clknet_leaf_6_wb_clk_i),
    .Q(\as2650.psu[4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _9390_ (.D(_0283_),
    .CLK(clknet_leaf_5_wb_clk_i),
    .Q(\as2650.psu[3] ));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _9432_ (.I(net46),
    .Z(net14));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _9433_ (.I(net46),
    .Z(net15));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _9434_ (.I(net47),
    .Z(net16));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _9435_ (.I(net47),
    .Z(net17));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _9436_ (.I(net46),
    .Z(net18));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _9437_ (.I(net47),
    .Z(net11));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _9438_ (.I(net46),
    .Z(net12));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_0_wb_clk_i (.I(wb_clk_i),
    .Z(clknet_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8 clkbuf_3_0_0_wb_clk_i (.I(clknet_0_wb_clk_i),
    .Z(clknet_3_0_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8 clkbuf_3_1_0_wb_clk_i (.I(clknet_0_wb_clk_i),
    .Z(clknet_3_1_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8 clkbuf_3_2_0_wb_clk_i (.I(clknet_0_wb_clk_i),
    .Z(clknet_3_2_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8 clkbuf_3_3_0_wb_clk_i (.I(clknet_0_wb_clk_i),
    .Z(clknet_3_3_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8 clkbuf_3_4_0_wb_clk_i (.I(clknet_0_wb_clk_i),
    .Z(clknet_3_4_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8 clkbuf_3_5_0_wb_clk_i (.I(clknet_0_wb_clk_i),
    .Z(clknet_3_5_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8 clkbuf_3_6_0_wb_clk_i (.I(clknet_0_wb_clk_i),
    .Z(clknet_3_6_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8 clkbuf_3_7_0_wb_clk_i (.I(clknet_0_wb_clk_i),
    .Z(clknet_3_7_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_11_wb_clk_i (.I(clknet_3_2_0_wb_clk_i),
    .Z(clknet_leaf_11_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_12_wb_clk_i (.I(clknet_3_2_0_wb_clk_i),
    .Z(clknet_leaf_12_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_14_wb_clk_i (.I(clknet_3_2_0_wb_clk_i),
    .Z(clknet_leaf_14_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_15_wb_clk_i (.I(clknet_3_2_0_wb_clk_i),
    .Z(clknet_leaf_15_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_16_wb_clk_i (.I(clknet_3_3_0_wb_clk_i),
    .Z(clknet_leaf_16_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_18_wb_clk_i (.I(clknet_3_3_0_wb_clk_i),
    .Z(clknet_leaf_18_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_1_wb_clk_i (.I(clknet_3_0_0_wb_clk_i),
    .Z(clknet_leaf_1_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_20_wb_clk_i (.I(clknet_3_3_0_wb_clk_i),
    .Z(clknet_leaf_20_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_23_wb_clk_i (.I(clknet_3_3_0_wb_clk_i),
    .Z(clknet_leaf_23_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_24_wb_clk_i (.I(clknet_3_6_0_wb_clk_i),
    .Z(clknet_leaf_24_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_25_wb_clk_i (.I(clknet_3_6_0_wb_clk_i),
    .Z(clknet_leaf_25_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_26_wb_clk_i (.I(clknet_opt_1_0_wb_clk_i),
    .Z(clknet_leaf_26_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_27_wb_clk_i (.I(clknet_3_6_0_wb_clk_i),
    .Z(clknet_leaf_27_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_28_wb_clk_i (.I(clknet_3_6_0_wb_clk_i),
    .Z(clknet_leaf_28_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_29_wb_clk_i (.I(clknet_3_6_0_wb_clk_i),
    .Z(clknet_leaf_29_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_2_wb_clk_i (.I(clknet_3_0_0_wb_clk_i),
    .Z(clknet_leaf_2_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_30_wb_clk_i (.I(clknet_3_6_0_wb_clk_i),
    .Z(clknet_leaf_30_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_31_wb_clk_i (.I(clknet_3_6_0_wb_clk_i),
    .Z(clknet_leaf_31_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_36_wb_clk_i (.I(clknet_3_7_0_wb_clk_i),
    .Z(clknet_leaf_36_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_37_wb_clk_i (.I(clknet_3_7_0_wb_clk_i),
    .Z(clknet_leaf_37_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_38_wb_clk_i (.I(clknet_3_7_0_wb_clk_i),
    .Z(clknet_leaf_38_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_39_wb_clk_i (.I(clknet_3_7_0_wb_clk_i),
    .Z(clknet_leaf_39_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_3_wb_clk_i (.I(clknet_3_2_0_wb_clk_i),
    .Z(clknet_leaf_3_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_40_wb_clk_i (.I(clknet_3_7_0_wb_clk_i),
    .Z(clknet_leaf_40_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_41_wb_clk_i (.I(clknet_3_7_0_wb_clk_i),
    .Z(clknet_leaf_41_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_42_wb_clk_i (.I(clknet_3_7_0_wb_clk_i),
    .Z(clknet_leaf_42_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_44_wb_clk_i (.I(clknet_3_5_0_wb_clk_i),
    .Z(clknet_leaf_44_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_45_wb_clk_i (.I(clknet_3_5_0_wb_clk_i),
    .Z(clknet_leaf_45_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_46_wb_clk_i (.I(clknet_3_4_0_wb_clk_i),
    .Z(clknet_leaf_46_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_47_wb_clk_i (.I(clknet_3_5_0_wb_clk_i),
    .Z(clknet_leaf_47_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_48_wb_clk_i (.I(clknet_3_5_0_wb_clk_i),
    .Z(clknet_leaf_48_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_49_wb_clk_i (.I(clknet_3_5_0_wb_clk_i),
    .Z(clknet_leaf_49_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_50_wb_clk_i (.I(clknet_3_5_0_wb_clk_i),
    .Z(clknet_leaf_50_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_51_wb_clk_i (.I(clknet_3_7_0_wb_clk_i),
    .Z(clknet_leaf_51_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_52_wb_clk_i (.I(clknet_3_5_0_wb_clk_i),
    .Z(clknet_leaf_52_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_53_wb_clk_i (.I(clknet_3_5_0_wb_clk_i),
    .Z(clknet_leaf_53_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_54_wb_clk_i (.I(clknet_3_5_0_wb_clk_i),
    .Z(clknet_leaf_54_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_55_wb_clk_i (.I(clknet_3_5_0_wb_clk_i),
    .Z(clknet_leaf_55_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_56_wb_clk_i (.I(clknet_3_5_0_wb_clk_i),
    .Z(clknet_leaf_56_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_57_wb_clk_i (.I(clknet_3_5_0_wb_clk_i),
    .Z(clknet_leaf_57_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_58_wb_clk_i (.I(clknet_3_5_0_wb_clk_i),
    .Z(clknet_leaf_58_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_59_wb_clk_i (.I(clknet_3_5_0_wb_clk_i),
    .Z(clknet_leaf_59_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_5_wb_clk_i (.I(clknet_3_1_0_wb_clk_i),
    .Z(clknet_leaf_5_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_60_wb_clk_i (.I(clknet_3_5_0_wb_clk_i),
    .Z(clknet_leaf_60_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_61_wb_clk_i (.I(clknet_3_5_0_wb_clk_i),
    .Z(clknet_leaf_61_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_62_wb_clk_i (.I(clknet_3_4_0_wb_clk_i),
    .Z(clknet_leaf_62_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_63_wb_clk_i (.I(clknet_3_4_0_wb_clk_i),
    .Z(clknet_leaf_63_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_64_wb_clk_i (.I(clknet_3_4_0_wb_clk_i),
    .Z(clknet_leaf_64_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_65_wb_clk_i (.I(clknet_3_4_0_wb_clk_i),
    .Z(clknet_leaf_65_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_66_wb_clk_i (.I(clknet_3_4_0_wb_clk_i),
    .Z(clknet_leaf_66_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_67_wb_clk_i (.I(clknet_3_4_0_wb_clk_i),
    .Z(clknet_leaf_67_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_68_wb_clk_i (.I(clknet_3_4_0_wb_clk_i),
    .Z(clknet_leaf_68_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_69_wb_clk_i (.I(clknet_3_4_0_wb_clk_i),
    .Z(clknet_leaf_69_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_6_wb_clk_i (.I(clknet_3_1_0_wb_clk_i),
    .Z(clknet_leaf_6_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_71_wb_clk_i (.I(clknet_3_4_0_wb_clk_i),
    .Z(clknet_leaf_71_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_73_wb_clk_i (.I(clknet_3_1_0_wb_clk_i),
    .Z(clknet_leaf_73_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_74_wb_clk_i (.I(clknet_3_1_0_wb_clk_i),
    .Z(clknet_leaf_74_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_75_wb_clk_i (.I(clknet_3_1_0_wb_clk_i),
    .Z(clknet_leaf_75_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_76_wb_clk_i (.I(clknet_3_1_0_wb_clk_i),
    .Z(clknet_leaf_76_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_77_wb_clk_i (.I(clknet_3_1_0_wb_clk_i),
    .Z(clknet_leaf_77_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_80_wb_clk_i (.I(clknet_3_0_0_wb_clk_i),
    .Z(clknet_leaf_80_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_8_wb_clk_i (.I(clknet_3_3_0_wb_clk_i),
    .Z(clknet_leaf_8_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_9_wb_clk_i (.I(clknet_3_3_0_wb_clk_i),
    .Z(clknet_leaf_9_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_opt_1_0_wb_clk_i (.I(clknet_3_6_0_wb_clk_i),
    .Z(clknet_opt_1_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 fanout46 (.I(net48),
    .Z(net46));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout47 (.I(net48),
    .Z(net47));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout48 (.I(net49),
    .Z(net48));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout49 (.I(net50),
    .Z(net49));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout50 (.I(net13),
    .Z(net50));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 fanout51 (.I(net25),
    .Z(net51));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 fanout52 (.I(net40),
    .Z(net52));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 fanout53 (.I(net38),
    .Z(net53));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 fanout54 (.I(net35),
    .Z(net54));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 input1 (.I(io_in[10]),
    .Z(net1));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 input10 (.I(io_in[9]),
    .Z(net10));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 input2 (.I(io_in[11]),
    .Z(net2));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input3 (.I(io_in[12]),
    .Z(net3));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 input4 (.I(io_in[13]),
    .Z(net4));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input5 (.I(io_in[33]),
    .Z(net5));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 input6 (.I(io_in[5]),
    .Z(net6));
 gf180mcu_fd_sc_mcu7t5v0__dlyd_1 input7 (.I(io_in[6]),
    .Z(net7));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 input8 (.I(io_in[7]),
    .Z(net8));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 input9 (.I(io_in[8]),
    .Z(net9));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output11 (.I(net11),
    .Z(io_oeb[10]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output12 (.I(net12),
    .Z(io_oeb[11]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output13 (.I(net50),
    .Z(io_oeb[12]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output14 (.I(net14),
    .Z(io_oeb[5]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output15 (.I(net15),
    .Z(io_oeb[6]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output16 (.I(net16),
    .Z(io_oeb[7]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output17 (.I(net17),
    .Z(io_oeb[8]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output18 (.I(net18),
    .Z(io_oeb[9]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output19 (.I(net19),
    .Z(io_out[10]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output20 (.I(net20),
    .Z(io_out[11]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output21 (.I(net21),
    .Z(io_out[12]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output22 (.I(net22),
    .Z(io_out[14]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output23 (.I(net23),
    .Z(io_out[15]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output24 (.I(net24),
    .Z(io_out[16]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output25 (.I(net25),
    .Z(io_out[17]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output26 (.I(net26),
    .Z(io_out[18]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output27 (.I(net27),
    .Z(io_out[19]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output28 (.I(net28),
    .Z(io_out[20]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output29 (.I(net29),
    .Z(io_out[21]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output30 (.I(net30),
    .Z(io_out[22]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output31 (.I(net31),
    .Z(io_out[23]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output32 (.I(net32),
    .Z(io_out[24]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output33 (.I(net33),
    .Z(io_out[25]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output34 (.I(net34),
    .Z(io_out[26]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output35 (.I(net35),
    .Z(io_out[27]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output36 (.I(net36),
    .Z(io_out[28]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output37 (.I(net37),
    .Z(io_out[29]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output38 (.I(net38),
    .Z(io_out[30]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output39 (.I(net39),
    .Z(io_out[31]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output40 (.I(net40),
    .Z(io_out[32]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output41 (.I(net41),
    .Z(io_out[5]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output42 (.I(net42),
    .Z(io_out[6]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output43 (.I(net43),
    .Z(io_out[7]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output44 (.I(net44),
    .Z(io_out[8]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output45 (.I(net45),
    .Z(io_out[9]));
 gf180mcu_fd_sc_mcu7t5v0__tiel wrapped_as2650_55 (.ZN(net55));
 gf180mcu_fd_sc_mcu7t5v0__tiel wrapped_as2650_56 (.ZN(net56));
 gf180mcu_fd_sc_mcu7t5v0__tiel wrapped_as2650_57 (.ZN(net57));
 gf180mcu_fd_sc_mcu7t5v0__tiel wrapped_as2650_58 (.ZN(net58));
 gf180mcu_fd_sc_mcu7t5v0__tiel wrapped_as2650_59 (.ZN(net59));
 gf180mcu_fd_sc_mcu7t5v0__tiel wrapped_as2650_60 (.ZN(net60));
 gf180mcu_fd_sc_mcu7t5v0__tiel wrapped_as2650_61 (.ZN(net61));
 gf180mcu_fd_sc_mcu7t5v0__tiel wrapped_as2650_62 (.ZN(net62));
 gf180mcu_fd_sc_mcu7t5v0__tiel wrapped_as2650_63 (.ZN(net63));
 gf180mcu_fd_sc_mcu7t5v0__tiel wrapped_as2650_64 (.ZN(net64));
 gf180mcu_fd_sc_mcu7t5v0__tiel wrapped_as2650_65 (.ZN(net65));
 gf180mcu_fd_sc_mcu7t5v0__tiel wrapped_as2650_66 (.ZN(net66));
 gf180mcu_fd_sc_mcu7t5v0__tiel wrapped_as2650_67 (.ZN(net67));
 gf180mcu_fd_sc_mcu7t5v0__tiel wrapped_as2650_68 (.ZN(net68));
 gf180mcu_fd_sc_mcu7t5v0__tiel wrapped_as2650_69 (.ZN(net69));
 gf180mcu_fd_sc_mcu7t5v0__tiel wrapped_as2650_70 (.ZN(net70));
 gf180mcu_fd_sc_mcu7t5v0__tiel wrapped_as2650_71 (.ZN(net71));
 gf180mcu_fd_sc_mcu7t5v0__tiel wrapped_as2650_72 (.ZN(net72));
 gf180mcu_fd_sc_mcu7t5v0__tiel wrapped_as2650_73 (.ZN(net73));
 gf180mcu_fd_sc_mcu7t5v0__tiel wrapped_as2650_74 (.ZN(net74));
 gf180mcu_fd_sc_mcu7t5v0__tiel wrapped_as2650_75 (.ZN(net75));
 gf180mcu_fd_sc_mcu7t5v0__tiel wrapped_as2650_76 (.ZN(net76));
 gf180mcu_fd_sc_mcu7t5v0__tiel wrapped_as2650_77 (.ZN(net77));
 gf180mcu_fd_sc_mcu7t5v0__tiel wrapped_as2650_78 (.ZN(net78));
 gf180mcu_fd_sc_mcu7t5v0__tiel wrapped_as2650_79 (.ZN(net79));
 gf180mcu_fd_sc_mcu7t5v0__tiel wrapped_as2650_80 (.ZN(net80));
 gf180mcu_fd_sc_mcu7t5v0__tiel wrapped_as2650_81 (.ZN(net81));
 gf180mcu_fd_sc_mcu7t5v0__tiel wrapped_as2650_82 (.ZN(net82));
 gf180mcu_fd_sc_mcu7t5v0__tiel wrapped_as2650_83 (.ZN(net83));
 gf180mcu_fd_sc_mcu7t5v0__tiel wrapped_as2650_84 (.ZN(net84));
 gf180mcu_fd_sc_mcu7t5v0__tieh wrapped_as2650_85 (.Z(net85));
 gf180mcu_fd_sc_mcu7t5v0__tieh wrapped_as2650_86 (.Z(net86));
 gf180mcu_fd_sc_mcu7t5v0__tieh wrapped_as2650_87 (.Z(net87));
 gf180mcu_fd_sc_mcu7t5v0__tieh wrapped_as2650_88 (.Z(net88));
 gf180mcu_fd_sc_mcu7t5v0__tieh wrapped_as2650_89 (.Z(net89));
 gf180mcu_fd_sc_mcu7t5v0__tieh wrapped_as2650_90 (.Z(net90));
 gf180mcu_fd_sc_mcu7t5v0__tieh wrapped_as2650_91 (.Z(net91));
 gf180mcu_fd_sc_mcu7t5v0__tieh wrapped_as2650_92 (.Z(net92));
 gf180mcu_fd_sc_mcu7t5v0__tieh wrapped_as2650_93 (.Z(net93));
 gf180mcu_fd_sc_mcu7t5v0__tieh wrapped_as2650_94 (.Z(net94));
 gf180mcu_fd_sc_mcu7t5v0__tieh wrapped_as2650_95 (.Z(net95));
 assign io_oeb[0] = net85;
 assign io_oeb[13] = net90;
 assign io_oeb[14] = net55;
 assign io_oeb[15] = net56;
 assign io_oeb[16] = net57;
 assign io_oeb[17] = net58;
 assign io_oeb[18] = net59;
 assign io_oeb[19] = net60;
 assign io_oeb[1] = net86;
 assign io_oeb[20] = net61;
 assign io_oeb[21] = net62;
 assign io_oeb[22] = net63;
 assign io_oeb[23] = net64;
 assign io_oeb[24] = net65;
 assign io_oeb[25] = net66;
 assign io_oeb[26] = net67;
 assign io_oeb[27] = net68;
 assign io_oeb[28] = net69;
 assign io_oeb[29] = net70;
 assign io_oeb[2] = net87;
 assign io_oeb[30] = net71;
 assign io_oeb[31] = net72;
 assign io_oeb[32] = net73;
 assign io_oeb[33] = net91;
 assign io_oeb[34] = net92;
 assign io_oeb[35] = net93;
 assign io_oeb[36] = net94;
 assign io_oeb[37] = net95;
 assign io_oeb[3] = net88;
 assign io_oeb[4] = net89;
 assign io_out[0] = net74;
 assign io_out[13] = net79;
 assign io_out[1] = net75;
 assign io_out[2] = net76;
 assign io_out[33] = net80;
 assign io_out[34] = net81;
 assign io_out[35] = net82;
 assign io_out[36] = net83;
 assign io_out[37] = net84;
 assign io_out[3] = net77;
 assign io_out[4] = net78;
endmodule

