// This is the unpowered netlist.
module ram_controller (CEN_all,
    GWEN_0,
    GWEN_1,
    GWEN_2,
    GWEN_3,
    GWEN_4,
    GWEN_5,
    GWEN_6,
    GWEN_7,
    WEb_raw,
    ram_enabled,
    rst,
    wb_clk_i,
    A_all,
    D_all,
    Q0,
    Q1,
    Q2,
    Q3,
    Q4,
    Q5,
    Q6,
    Q7,
    WEN_all,
    bus_in,
    bus_out,
    requested_addr);
 output CEN_all;
 output GWEN_0;
 output GWEN_1;
 output GWEN_2;
 output GWEN_3;
 output GWEN_4;
 output GWEN_5;
 output GWEN_6;
 output GWEN_7;
 input WEb_raw;
 input ram_enabled;
 input rst;
 input wb_clk_i;
 output [8:0] A_all;
 output [7:0] D_all;
 input [7:0] Q0;
 input [7:0] Q1;
 input [7:0] Q2;
 input [7:0] Q3;
 input [7:0] Q4;
 input [7:0] Q5;
 input [7:0] Q6;
 input [7:0] Q7;
 output [7:0] WEN_all;
 input [7:0] bus_in;
 output [7:0] bus_out;
 input [15:0] requested_addr;

 wire net126;
 wire net127;
 wire net128;
 wire net129;
 wire net130;
 wire net131;
 wire net132;
 wire net133;
 wire _000_;
 wire _001_;
 wire _002_;
 wire _003_;
 wire _004_;
 wire _005_;
 wire _006_;
 wire _007_;
 wire _008_;
 wire _009_;
 wire _010_;
 wire _011_;
 wire _012_;
 wire _013_;
 wire _014_;
 wire _015_;
 wire _016_;
 wire _017_;
 wire _018_;
 wire _019_;
 wire _020_;
 wire _021_;
 wire _022_;
 wire _023_;
 wire _024_;
 wire _025_;
 wire _026_;
 wire _027_;
 wire _028_;
 wire _029_;
 wire _030_;
 wire _031_;
 wire _032_;
 wire _033_;
 wire _034_;
 wire _035_;
 wire _036_;
 wire _037_;
 wire _038_;
 wire _039_;
 wire _040_;
 wire _041_;
 wire _042_;
 wire _043_;
 wire _044_;
 wire _045_;
 wire _046_;
 wire _047_;
 wire _048_;
 wire _049_;
 wire _050_;
 wire _051_;
 wire _052_;
 wire _053_;
 wire _054_;
 wire _055_;
 wire _056_;
 wire _057_;
 wire _058_;
 wire _059_;
 wire _060_;
 wire _061_;
 wire _062_;
 wire _063_;
 wire _064_;
 wire _065_;
 wire _066_;
 wire _067_;
 wire _068_;
 wire _069_;
 wire _070_;
 wire _071_;
 wire _072_;
 wire _073_;
 wire _074_;
 wire _075_;
 wire _076_;
 wire _077_;
 wire _078_;
 wire _079_;
 wire _080_;
 wire _081_;
 wire _082_;
 wire _083_;
 wire _084_;
 wire _085_;
 wire _086_;
 wire _087_;
 wire _088_;
 wire _089_;
 wire _090_;
 wire _091_;
 wire _092_;
 wire _093_;
 wire _094_;
 wire _095_;
 wire _096_;
 wire _097_;
 wire _098_;
 wire _099_;
 wire _100_;
 wire _101_;
 wire _102_;
 wire _103_;
 wire _104_;
 wire _105_;
 wire \aaaa[0] ;
 wire \aaaa[10] ;
 wire \aaaa[11] ;
 wire \aaaa[12] ;
 wire \aaaa[13] ;
 wire \aaaa[14] ;
 wire \aaaa[15] ;
 wire \aaaa[1] ;
 wire \aaaa[2] ;
 wire \aaaa[3] ;
 wire \aaaa[4] ;
 wire \aaaa[5] ;
 wire \aaaa[6] ;
 wire \aaaa[7] ;
 wire \aaaa[8] ;
 wire \aaaa[9] ;
 wire clknet_0_wb_clk_i;
 wire clknet_1_0__leaf_wb_clk_i;
 wire clknet_1_1__leaf_wb_clk_i;
 wire net1;
 wire net10;
 wire net100;
 wire net101;
 wire net102;
 wire net103;
 wire net104;
 wire net105;
 wire net106;
 wire net107;
 wire net108;
 wire net109;
 wire net11;
 wire net110;
 wire net111;
 wire net112;
 wire net113;
 wire net114;
 wire net115;
 wire net116;
 wire net117;
 wire net118;
 wire net119;
 wire net12;
 wire net120;
 wire net121;
 wire net122;
 wire net123;
 wire net124;
 wire net125;
 wire net13;
 wire net14;
 wire net15;
 wire net16;
 wire net17;
 wire net18;
 wire net19;
 wire net2;
 wire net20;
 wire net21;
 wire net22;
 wire net23;
 wire net24;
 wire net25;
 wire net26;
 wire net27;
 wire net28;
 wire net29;
 wire net3;
 wire net30;
 wire net31;
 wire net32;
 wire net33;
 wire net34;
 wire net35;
 wire net36;
 wire net37;
 wire net38;
 wire net39;
 wire net4;
 wire net40;
 wire net41;
 wire net42;
 wire net43;
 wire net44;
 wire net45;
 wire net46;
 wire net47;
 wire net48;
 wire net49;
 wire net5;
 wire net50;
 wire net51;
 wire net52;
 wire net53;
 wire net54;
 wire net55;
 wire net56;
 wire net57;
 wire net58;
 wire net59;
 wire net6;
 wire net60;
 wire net61;
 wire net62;
 wire net63;
 wire net64;
 wire net65;
 wire net66;
 wire net67;
 wire net68;
 wire net69;
 wire net7;
 wire net70;
 wire net71;
 wire net72;
 wire net73;
 wire net74;
 wire net75;
 wire net76;
 wire net77;
 wire net78;
 wire net79;
 wire net8;
 wire net80;
 wire net81;
 wire net82;
 wire net83;
 wire net84;
 wire net85;
 wire net86;
 wire net87;
 wire net88;
 wire net89;
 wire net9;
 wire net90;
 wire net91;
 wire net92;
 wire net93;
 wire net94;
 wire net95;
 wire net96;
 wire net97;
 wire net98;
 wire net99;

 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__108__A4 (.I(net52));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__109__A1 (.I(_068_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__110__B2 (.I(_076_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__111__I (.I(net5));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__112__B2 (.I(net45));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__112__C1 (.I(net61));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__113__A4 (.I(net13));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__115__A2 (.I(net37));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__116__A4 (.I(net53));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__117__A1 (.I(_079_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__118__B2 (.I(_083_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__119__I (.I(net6));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__120__B2 (.I(net46));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__120__C1 (.I(net62));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__121__A4 (.I(net14));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__123__A2 (.I(net38));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__124__A4 (.I(net54));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__125__A1 (.I(_086_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__126__B2 (.I(_090_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__127__I (.I(net7));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__128__B2 (.I(net47));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__128__C1 (.I(net63));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__129__A4 (.I(net15));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__131__A2 (.I(net39));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__132__A4 (.I(net55));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__134__B2 (.I(_097_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__135__I (.I(net8));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__136__B1 (.I(_026_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__136__B2 (.I(net48));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__136__C1 (.I(net64));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__137__A4 (.I(net16));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__138__A2 (.I(net32));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__138__A3 (.I(_020_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__139__A2 (.I(net40));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__140__A4 (.I(net56));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__142__A2 (.I(_009_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__142__B1 (.I(_099_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__142__B2 (.I(_104_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__144__A1 (.I(net74));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__145__A1 (.I(net65));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__146__I (.I(_001_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__147__I (.I(\aaaa[1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__149__I (.I(\aaaa[0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__151__I (.I(\aaaa[2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__154__I (.I(_009_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__159__I (.I(\aaaa[2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__162__I (.I(_001_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__163__A4 (.I(_017_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__167__A1 (.I(\aaaa[1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__167__A2 (.I(\aaaa[0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__168__I (.I(_020_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__169__A2 (.I(_017_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__173__A2 (.I(_017_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__176__I (.I(_026_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__180__A4 (.I(_017_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__181__A2 (.I(_020_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__184__I (.I(net1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__185__B2 (.I(net41));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__185__C1 (.I(net57));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__188__A4 (.I(net9));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__191__A2 (.I(net33));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__192__A4 (.I(net49));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__194__B2 (.I(_041_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__195__I (.I(net2));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__196__B2 (.I(net42));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__196__C1 (.I(net58));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__197__A4 (.I(net10));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__199__A2 (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__200__A4 (.I(net50));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__202__B2 (.I(_048_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__203__I (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__204__B2 (.I(net43));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__204__C1 (.I(net59));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__206__A4 (.I(net11));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__210__A2 (.I(net35));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__212__A4 (.I(net51));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__214__B2 (.I(_059_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__215__I (.I(net4));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__216__I (.I(_009_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__218__I (.I(_026_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__220__B2 (.I(net44));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__220__C1 (.I(net60));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__223__A4 (.I(net12));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__224__I (.I(_020_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__227__A2 (.I(net36));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__228__CLK (.I(clknet_1_1__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__228__D (.I(net75));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__229__CLK (.I(clknet_1_1__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__229__D (.I(net82));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__230__CLK (.I(clknet_1_1__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__230__D (.I(net83));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__231__CLK (.I(clknet_1_0__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__232__CLK (.I(clknet_1_0__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__233__CLK (.I(clknet_1_0__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__234__CLK (.I(clknet_1_0__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__235__CLK (.I(clknet_1_0__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__236__CLK (.I(clknet_1_0__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__237__CLK (.I(clknet_1_0__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__238__CLK (.I(clknet_1_1__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__239__CLK (.I(clknet_1_1__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__240__CLK (.I(clknet_1_1__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__241__CLK (.I(clknet_1_1__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__242__CLK (.I(clknet_1_1__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__243__CLK (.I(clknet_1_1__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__261__I (.I(net91));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__262__I (.I(net66));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__263__I (.I(net67));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__264__I (.I(net68));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__265__I (.I(net69));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__266__I (.I(net70));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__267__I (.I(net71));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__268__I (.I(net72));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__269__I (.I(net73));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_0_wb_clk_i_I (.I(wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_1_0__f_wb_clk_i_I (.I(clknet_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_1_1__f_wb_clk_i_I (.I(clknet_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input10_I (.I(Q1[1]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input11_I (.I(Q1[2]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input12_I (.I(Q1[3]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input13_I (.I(Q1[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input14_I (.I(Q1[5]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input15_I (.I(Q1[6]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input16_I (.I(Q1[7]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input17_I (.I(Q2[0]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input18_I (.I(Q2[1]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input19_I (.I(Q2[2]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input1_I (.I(Q0[0]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input20_I (.I(Q2[3]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input21_I (.I(Q2[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input22_I (.I(Q2[5]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input23_I (.I(Q2[6]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input24_I (.I(Q2[7]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input25_I (.I(Q3[0]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input26_I (.I(Q3[1]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input27_I (.I(Q3[2]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input28_I (.I(Q3[3]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input29_I (.I(Q3[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input2_I (.I(Q0[1]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input30_I (.I(Q3[5]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input31_I (.I(Q3[6]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input32_I (.I(Q3[7]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input33_I (.I(Q4[0]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input34_I (.I(Q4[1]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input35_I (.I(Q4[2]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input36_I (.I(Q4[3]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input37_I (.I(Q4[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input38_I (.I(Q4[5]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input39_I (.I(Q4[6]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input3_I (.I(Q0[2]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input40_I (.I(Q4[7]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input41_I (.I(Q5[0]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input42_I (.I(Q5[1]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input43_I (.I(Q5[2]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input44_I (.I(Q5[3]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input45_I (.I(Q5[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input46_I (.I(Q5[5]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input47_I (.I(Q5[6]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input48_I (.I(Q5[7]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input49_I (.I(Q6[0]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input4_I (.I(Q0[3]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input50_I (.I(Q6[1]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input51_I (.I(Q6[2]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input52_I (.I(Q6[3]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input53_I (.I(Q6[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input54_I (.I(Q6[5]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input55_I (.I(Q6[6]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input56_I (.I(Q6[7]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input57_I (.I(Q7[0]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input58_I (.I(Q7[1]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input59_I (.I(Q7[2]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input5_I (.I(Q0[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input60_I (.I(Q7[3]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input61_I (.I(Q7[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input62_I (.I(Q7[5]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input63_I (.I(Q7[6]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input64_I (.I(Q7[7]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input65_I (.I(WEb_raw));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input66_I (.I(bus_in[0]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input67_I (.I(bus_in[1]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input68_I (.I(bus_in[2]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input69_I (.I(bus_in[3]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input6_I (.I(Q0[5]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input70_I (.I(bus_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input71_I (.I(bus_in[5]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input72_I (.I(bus_in[6]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input73_I (.I(bus_in[7]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input74_I (.I(ram_enabled));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input75_I (.I(requested_addr[0]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input76_I (.I(requested_addr[10]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input77_I (.I(requested_addr[11]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input78_I (.I(requested_addr[12]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input79_I (.I(requested_addr[13]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input7_I (.I(Q0[6]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input80_I (.I(requested_addr[14]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input81_I (.I(requested_addr[15]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input82_I (.I(requested_addr[1]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input83_I (.I(requested_addr[2]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input84_I (.I(requested_addr[3]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input85_I (.I(requested_addr[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input86_I (.I(requested_addr[5]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input87_I (.I(requested_addr[6]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input88_I (.I(requested_addr[7]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input89_I (.I(requested_addr[8]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input8_I (.I(Q0[7]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input90_I (.I(requested_addr[9]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input91_I (.I(rst));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input9_I (.I(Q1[0]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output100_I (.I(net100));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output110_I (.I(net110));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output111_I (.I(net111));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output112_I (.I(net112));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output113_I (.I(net113));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output114_I (.I(net114));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output115_I (.I(net115));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output116_I (.I(net116));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output117_I (.I(net117));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output118_I (.I(net118));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output119_I (.I(net119));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output120_I (.I(net120));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output121_I (.I(net121));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output122_I (.I(net122));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output123_I (.I(net123));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output124_I (.I(net124));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output125_I (.I(net125));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output92_I (.I(net92));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output93_I (.I(net93));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output94_I (.I(net94));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output95_I (.I(net95));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output96_I (.I(net96));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output97_I (.I(net97));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output98_I (.I(net98));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output99_I (.I(net99));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_0_100 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_0_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_0_1019 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_0_1022 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_0_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_0_1049 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_0_1053 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_0_1082 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_0_1096 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_0_1112 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_0_1130 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_0_1146 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_0_1164 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_0_1180 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_0_1189 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_0_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_0_120 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_0_1208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_0_1212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_0_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_0_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_0_1226 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_0_124 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_0_1242 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_0_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_0_1253 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_0_1257 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_0_126 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_0_1260 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_0_1276 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_0_1285 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_0_1289 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_0_1291 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_0_1294 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_0_1302 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_0_1306 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_0_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_0_131 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_0_1317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_0_1325 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_0_1328 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_0_1336 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_0_1340 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_0_1349 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_0_135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_0_1357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_0_1359 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_0_1362 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_0_1370 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_0_1372 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_0_138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_0_1381 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_0_1389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_0_1393 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_0_1396 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_0_1404 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_0_1413 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_0_1421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_0_1425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_0_1427 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_0_1430 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_0_1434 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_0_1436 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_0_1445 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_0_1461 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_0_1464 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_0_1468 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_0_1477 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_0_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_0_1495 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_0_1498 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_0_1500 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_0_1509 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_0_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_0_1527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_0_1532 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_0_1534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_0_154 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_0_1541 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_0_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_0_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_0_1566 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_0_1573 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_0_158 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_0_1589 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_0_1593 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_0_1595 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_0_1606 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_0_1610 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_0_1618 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_0_1622 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_0_163 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_0_1650 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_0_1656 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_0_167 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_0_1674 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_0_1682 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_0_1686 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_0_169 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_0_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_0_1742 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_0_1746 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_0_1750 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_0_1754 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_0_1758 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_0_1765 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_0_1767 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_0_1770 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_0_1774 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_0_1778 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_0_1782 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_0_1812 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_0_1831 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_0_1835 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_0_1844 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_0_1848 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_0_1852 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_0_1866 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_0_1879 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_0_188 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_0_1883 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_0_1893 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_0_190 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_0_1901 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_0_1903 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_0_1906 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_0_1912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_0_1916 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_0_1918 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_0_1925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_0_1933 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_0_1937 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_0_1940 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_0_1944 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_0_195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_0_1967 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_0_1971 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_0_1974 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_0_1978 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_0_1980 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_0_1989 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_0_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_0_2005 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_0_2008 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_0_2012 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_0_2021 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_0_203 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_0_2037 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_0_2039 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_0_2042 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_0_2044 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_0_2053 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_0_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_0_2069 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_0_2071 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_0_2076 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_0_2078 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_0_2085 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_0_2101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_0_2105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_0_2110 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_0_2117 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_0_2133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_0_2137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_0_2139 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_0_2150 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_0_2166 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_0_2184 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_0_2200 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_0_2218 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_0_222 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_0_2234 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_0_2252 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_0_2268 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_0_227 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_0_2277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_0_2280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_0_2296 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_0_2300 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_0_2309 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_0_2311 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_0_2314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_0_2330 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_0_2332 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_0_2341 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_0_2345 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_0_2348 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_0_235 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_0_2364 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_0_237 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_0_2375 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_0_2379 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_0_2382 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_0_2390 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_0_2394 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_0_2396 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_0_240 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_0_2407 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_0_2411 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_0_2413 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_0_2416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_0_2424 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_0_2428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_0_2439 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_0_2447 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_0_2450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_0_2458 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_0_2460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_0_2471 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_0_2479 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_0_248 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_0_2481 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_0_2484 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_0_2492 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_0_2503 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_0_2511 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_0_2515 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_0_2518 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_0_252 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_0_2522 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_0_2524 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_0_2535 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_0_254 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_0_2543 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_0_2547 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_0_2549 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_0_2552 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_0_2556 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_0_2567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_0_2583 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_0_2586 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_0_2588 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_0_259 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_0_2599 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_0_2615 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_0_2617 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_0_2620 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_0_267 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_0_271 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_0_274 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_0_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_0_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_0_291 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_0_299 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_0_303 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_0_305 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_0_308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_0_316 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_0_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_0_323 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_0_339 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_0_342 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_0_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_0_36 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_0_376 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_0_380 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_0_410 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_0_414 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_0_441 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_0_444 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_0_446 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_0_473 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_0_475 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_0_478 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_0_505 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_0_509 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_0_538 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_0_542 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_0_572 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_0_576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_0_606 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_0_610 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_0_640 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_0_644 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_0_674 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_0_678 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_0_682 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_0_686 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_0_695 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_0_711 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_0_713 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_0_716 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_0_724 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_0_726 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_0_729 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_0_745 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_0_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_0_750 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_0_758 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_0_761 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_0_777 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_0_779 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_0_790 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_0_806 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_0_814 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_0_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_0_822 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_0_852 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_0_856 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_0_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_0_890 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_0_920 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_0_924 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_0_954 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_0_958 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_0_985 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_0_988 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_0_990 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_10_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_10_1011 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_10_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_10_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_10_1081 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_10_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_10_1151 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_10_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_10_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_10_1227 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_10_1291 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_10_1297 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_10_1361 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_10_1367 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_10_1431 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_10_1437 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_10_1501 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_10_1507 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_10_1571 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_10_1577 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_10_1641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_10_1647 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_10_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_10_1711 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_10_1717 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_10_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_10_1781 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_10_1787 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_10_1851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_10_1857 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_10_1921 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_10_1927 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_10_1991 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_10_1997 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_10_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_10_2061 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_10_2067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_10_2131 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_10_2137 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_10_2201 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_10_2207 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_10_2271 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_10_2277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_10_2341 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_10_2347 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_10_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_10_2411 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_10_2417 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_10_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_10_2481 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_10_2487 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_10_2551 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_10_2557 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_10_2621 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_10_2627 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_10_2643 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_10_2651 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_10_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_10_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_10_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_10_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_10_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_10_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_10_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_10_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_10_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_10_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_10_591 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_10_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_10_661 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_10_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_10_731 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_10_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_10_801 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_10_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_10_871 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_10_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_10_941 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_10_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_11_1046 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_11_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_11_1116 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_11_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_11_1186 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_11_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_11_1256 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_11_1262 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_11_1326 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_11_1332 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_11_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_11_1396 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_11_1402 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_11_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_11_1466 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_11_1472 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_11_1536 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_11_1542 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_11_1606 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_11_1612 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_11_1676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_11_1682 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_11_1746 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_11_1752 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_11_1816 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_11_1822 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_11_1886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_11_1892 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_11_1956 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_11_1962 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_11_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_11_2026 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_11_2032 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_11_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_11_2096 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_11_2102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_11_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_11_2166 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_11_2172 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_11_2236 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_11_2242 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_11_2306 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_11_2312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_11_2376 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_11_2382 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_11_2446 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_11_2452 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_11_2516 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_11_2522 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_11_2586 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_11_2592 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_11_2624 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_11_2640 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_11_2648 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_11_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_11_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_11_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_11_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_11_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_11_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_11_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_11_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_11_556 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_11_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_11_626 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_11_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_11_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_11_696 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_11_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_11_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_11_766 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_11_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_11_836 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_11_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_11_906 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_11_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_11_976 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_11_982 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_12_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_12_1011 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_12_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_12_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_12_1081 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_12_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_12_1151 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_12_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_12_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_12_1227 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_12_1291 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_12_1297 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_12_1361 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_12_1367 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_12_1431 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_12_1437 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_12_1501 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_12_1507 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_12_1571 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_12_1577 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_12_1641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_12_1647 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_12_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_12_1711 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_12_1717 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_12_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_12_1781 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_12_1787 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_12_1851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_12_1857 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_12_1921 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_12_1927 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_12_1991 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_12_1997 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_12_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_12_2061 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_12_2067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_12_2131 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_12_2137 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_12_2201 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_12_2207 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_12_2271 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_12_2277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_12_2341 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_12_2347 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_12_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_12_2411 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_12_2417 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_12_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_12_2481 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_12_2487 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_12_2551 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_12_2557 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_12_2621 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_12_2627 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_12_2643 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_12_2651 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_12_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_12_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_12_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_12_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_12_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_12_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_12_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_12_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_12_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_12_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_12_591 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_12_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_12_661 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_12_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_12_731 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_12_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_12_801 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_12_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_12_871 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_12_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_12_941 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_12_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_13_1046 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_13_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_13_1116 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_13_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_13_1186 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_13_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_13_1256 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_13_1262 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_13_1326 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_13_1332 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_13_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_13_1396 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_13_1402 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_13_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_13_1466 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_13_1472 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_13_1536 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_13_1542 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_13_1606 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_13_1612 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_13_1676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_13_1682 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_13_1746 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_13_1752 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_13_1816 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_13_1822 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_13_1886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_13_1892 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_13_1956 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_13_1962 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_13_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_13_2026 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_13_2032 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_13_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_13_2096 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_13_2102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_13_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_13_2166 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_13_2172 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_13_2236 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_13_2242 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_13_2306 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_13_2312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_13_2376 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_13_2382 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_13_2446 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_13_2452 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_13_2516 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_13_2522 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_13_2586 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_13_2592 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_13_2624 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_13_2640 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_13_2648 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_13_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_13_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_13_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_13_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_13_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_13_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_13_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_13_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_13_556 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_13_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_13_626 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_13_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_13_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_13_696 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_13_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_13_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_13_766 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_13_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_13_836 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_13_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_13_906 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_13_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_13_976 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_13_982 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_14_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_14_1011 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_14_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_14_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_14_1081 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_14_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_14_1151 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_14_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_14_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_14_1227 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_14_1291 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_14_1297 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_14_1361 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_14_1367 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_14_1431 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_14_1437 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_14_1501 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_14_1507 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_14_1571 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_14_1577 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_14_1641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_14_1647 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_14_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_14_1711 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_14_1717 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_14_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_14_1781 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_14_1787 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_14_1851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_14_1857 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_14_1921 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_14_1927 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_14_1991 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_14_1997 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_14_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_14_2061 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_14_2067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_14_2131 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_14_2137 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_14_2201 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_14_2207 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_14_2271 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_14_2277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_14_2341 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_14_2347 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_14_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_14_2411 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_14_2417 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_14_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_14_2481 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_14_2487 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_14_2551 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_14_2557 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_14_2621 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_14_2627 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_14_2643 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_14_2651 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_14_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_14_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_14_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_14_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_14_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_14_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_14_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_14_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_14_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_14_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_14_591 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_14_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_14_661 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_14_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_14_731 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_14_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_14_801 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_14_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_14_871 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_14_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_14_941 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_14_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_15_1046 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_15_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_15_1116 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_15_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_15_1186 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_15_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_15_1256 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_15_1262 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_15_1326 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_15_1332 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_15_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_15_1396 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_15_1402 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_15_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_15_1466 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_15_1472 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_15_1536 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_15_1542 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_15_1606 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_15_1612 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_15_1676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_15_1682 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_15_1746 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_15_1752 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_15_1816 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_15_1822 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_15_1886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_15_1892 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_15_1956 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_15_1962 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_15_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_15_2026 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_15_2032 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_15_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_15_2096 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_15_2102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_15_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_15_2166 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_15_2172 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_15_2236 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_15_2242 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_15_2306 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_15_2312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_15_2376 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_15_2382 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_15_2446 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_15_2452 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_15_2516 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_15_2522 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_15_2586 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_15_2592 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_15_2624 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_15_2640 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_15_2648 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_15_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_15_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_15_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_15_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_15_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_15_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_15_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_15_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_15_556 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_15_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_15_626 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_15_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_15_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_15_696 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_15_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_15_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_15_766 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_15_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_15_836 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_15_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_15_906 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_15_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_15_976 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_15_982 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_16_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_16_1011 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_16_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_16_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_16_1081 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_16_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_16_1151 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_16_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_16_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_16_1227 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_16_1291 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_16_1297 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_16_1361 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_16_1367 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_16_1431 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_16_1437 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_16_1501 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_16_1507 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_16_1571 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_16_1577 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_16_1641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_16_1647 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_16_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_16_1711 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_16_1717 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_16_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_16_1781 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_16_1787 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_16_1851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_16_1857 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_16_1921 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_16_1927 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_16_1991 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_16_1997 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_16_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_16_2061 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_16_2067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_16_2131 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_16_2137 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_16_2201 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_16_2207 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_16_2271 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_16_2277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_16_2341 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_16_2347 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_16_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_16_2411 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_16_2417 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_16_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_16_2481 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_16_2487 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_16_2551 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_16_2557 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_16_2621 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_16_2627 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_16_2643 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_16_2651 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_16_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_16_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_16_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_16_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_16_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_16_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_16_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_16_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_16_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_16_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_16_591 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_16_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_16_661 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_16_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_16_731 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_16_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_16_801 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_16_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_16_871 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_16_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_16_941 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_16_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_17_1046 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_17_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_17_1116 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_17_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_17_1186 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_17_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_17_1256 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_17_1262 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_17_1326 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_17_1332 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_17_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_17_1396 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_17_1402 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_17_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_17_1466 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_17_1472 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_17_1536 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_17_1542 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_17_1606 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_17_1612 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_17_1676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_17_1682 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_17_1746 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_17_1752 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_17_1816 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_17_1822 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_17_1886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_17_1892 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_17_1956 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_17_1962 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_17_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_17_2026 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_17_2032 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_17_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_17_2096 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_17_2102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_17_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_17_2166 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_17_2172 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_17_2236 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_17_2242 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_17_2306 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_17_2312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_17_2376 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_17_2382 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_17_2446 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_17_2452 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_17_2516 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_17_2522 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_17_2586 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_17_2592 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_17_2624 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_17_2640 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_17_2648 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_17_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_17_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_17_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_17_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_17_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_17_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_17_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_17_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_17_556 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_17_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_17_626 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_17_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_17_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_17_696 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_17_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_17_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_17_766 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_17_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_17_836 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_17_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_17_906 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_17_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_17_976 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_17_982 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_18_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_18_1011 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_18_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_18_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_18_1081 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_18_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_18_1151 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_18_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_18_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_18_1227 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_18_1291 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_18_1297 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_18_1361 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_18_1367 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_18_1431 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_18_1437 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_18_1501 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_18_1507 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_18_1571 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_18_1577 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_18_1641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_18_1647 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_18_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_18_1711 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_18_1717 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_18_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_18_1781 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_18_1787 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_18_1851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_18_1857 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_18_1921 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_18_1927 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_18_1991 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_18_1997 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_18_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_18_2061 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_18_2067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_18_2131 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_18_2137 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_18_2201 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_18_2207 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_18_2271 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_18_2277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_18_2341 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_18_2347 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_18_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_18_2411 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_18_2417 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_18_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_18_2481 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_18_2487 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_18_2551 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_18_2557 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_18_2621 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_18_2627 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_18_2643 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_18_2651 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_18_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_18_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_18_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_18_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_18_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_18_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_18_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_18_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_18_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_18_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_18_591 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_18_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_18_661 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_18_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_18_731 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_18_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_18_801 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_18_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_18_871 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_18_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_18_941 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_18_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_19_1046 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_19_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_19_1116 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_19_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_19_1186 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_19_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_19_1256 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_19_1262 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_19_1326 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_19_1332 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_19_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_19_1396 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_19_1402 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_19_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_19_1466 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_19_1472 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_19_1536 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_19_1542 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_19_1606 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_19_1612 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_19_1676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_19_1682 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_19_1746 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_19_1752 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_19_1816 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_19_1822 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_19_1886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_19_1892 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_19_1956 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_19_1962 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_19_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_19_2026 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_19_2032 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_19_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_19_2096 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_19_2102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_19_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_19_2166 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_19_2172 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_19_2236 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_19_2242 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_19_2306 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_19_2312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_19_2376 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_19_2382 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_19_2446 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_19_2452 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_19_2516 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_19_2522 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_19_2586 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_19_2592 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_19_2624 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_19_2640 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_19_2648 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_19_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_19_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_19_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_19_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_19_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_19_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_19_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_19_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_19_556 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_19_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_19_626 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_19_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_19_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_19_696 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_19_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_19_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_19_766 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_19_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_19_836 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_19_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_19_906 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_19_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_19_976 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_19_982 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_1_100 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_1_1003 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_1_1011 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1_1015 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_1_1019 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_1_1035 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_1_1043 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1_1047 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1_1049 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_1_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_1_1068 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_1_1076 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1_1080 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_1_1084 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_1_1116 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_1_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_1_1186 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_1_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_1_1256 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_1_1262 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_1_132 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_1_1326 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_1_1332 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_1_1396 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_1_1402 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_1_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_1_1466 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_1_1472 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_1_1536 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_1_1542 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1_1606 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1_1612 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_1_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1_1729 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1_1733 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1_1737 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1_1739 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1_1815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1_1819 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1_1887 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1_1889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_1_1892 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_1_1900 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1_1904 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1_1914 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1_1918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1_1932 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_1_1936 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1_1944 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1_1955 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1_1957 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1_1973 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1_1983 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_1_1987 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_1_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_1_2019 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1_2027 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1_2029 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_1_2032 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_1_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_1_2096 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_1_2102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_1_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_1_2166 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_1_2172 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_1_2236 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_1_2242 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_1_2306 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_1_2312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_1_2376 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_1_2382 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_1_2446 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_1_2452 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_1_2516 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_1_2522 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_1_2586 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_1_2592 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_1_2624 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_1_2640 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_1_2648 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_1_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_1_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_1_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_1_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_1_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_1_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1_438 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1_440 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_1_443 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_1_459 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_1_467 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1_471 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_1_475 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_1_483 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1_487 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_1_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_1_556 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_1_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_1_594 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_1_610 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_1_618 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_1_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_1_648 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1_652 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1_654 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_1_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_1_663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1_697 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1_699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_1_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1_767 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1_769 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1_798 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_1_831 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1_839 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_1_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_1_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1_88 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_1_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_1_902 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_1_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1_96 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_1_976 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1_982 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1_984 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_1_987 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_20_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_20_1011 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_20_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_20_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_20_1081 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_20_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_20_1151 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_20_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_20_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_20_1227 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_20_1291 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_20_1297 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_20_1361 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_20_1367 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_20_1431 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_20_1437 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_20_1501 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_20_1507 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_20_1571 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_20_1577 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_20_1641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_20_1647 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_20_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_20_1711 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_20_1717 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_20_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_20_1781 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_20_1787 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_20_1851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_20_1857 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_20_1921 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_20_1927 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_20_1991 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_20_1997 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_20_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_20_2061 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_20_2067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_20_2131 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_20_2137 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_20_2201 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_20_2207 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_20_2271 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_20_2277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_20_2341 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_20_2347 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_20_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_20_2411 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_20_2417 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_20_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_20_2481 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_20_2487 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_20_2551 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_20_2557 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_20_2621 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_20_2627 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_20_2643 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_20_2651 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_20_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_20_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_20_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_20_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_20_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_20_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_20_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_20_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_20_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_20_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_20_591 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_20_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_20_661 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_20_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_20_731 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_20_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_20_801 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_20_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_20_871 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_20_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_20_941 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_20_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_21_1046 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_21_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_21_1116 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_21_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_21_1186 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_21_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_21_1256 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_21_1262 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_21_1326 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_21_1332 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_21_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_21_1396 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_21_1402 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_21_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_21_1466 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_21_1472 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_21_1536 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_21_1542 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_21_1606 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_21_1612 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_21_1676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_21_1682 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_21_1746 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_21_1752 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_21_1816 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_21_1822 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_21_1886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_21_1892 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_21_1956 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_21_1962 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_21_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_21_2026 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_21_2032 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_21_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_21_2096 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_21_2102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_21_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_21_2166 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_21_2172 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_21_2236 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_21_2242 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_21_2306 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_21_2312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_21_2376 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_21_2382 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_21_2446 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_21_2452 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_21_2516 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_21_2522 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_21_2586 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_21_2592 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_21_2624 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_21_2640 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_21_2648 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_21_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_21_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_21_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_21_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_21_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_21_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_21_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_21_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_21_556 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_21_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_21_626 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_21_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_21_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_21_696 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_21_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_21_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_21_766 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_21_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_21_836 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_21_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_21_906 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_21_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_21_976 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_21_982 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_22_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_22_1011 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_22_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_22_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_22_1081 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_22_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_22_1151 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_22_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_22_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_22_1227 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_22_1291 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_22_1297 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_22_1361 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_22_1367 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_22_1431 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_22_1437 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_22_1501 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_22_1507 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_22_1571 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_22_1577 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_22_1641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_22_1647 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_22_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_22_1711 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_22_1717 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_22_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_22_1781 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_22_1787 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_22_1851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_22_1857 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_22_1921 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_22_1927 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_22_1991 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_22_1997 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_22_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_22_2061 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_22_2067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_22_2131 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_22_2137 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_22_2201 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_22_2207 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_22_2271 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_22_2277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_22_2341 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_22_2347 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_22_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_22_2411 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_22_2417 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_22_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_22_2481 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_22_2487 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_22_2551 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_22_2557 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_22_2621 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_22_2627 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_22_2643 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_22_2651 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_22_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_22_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_22_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_22_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_22_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_22_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_22_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_22_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_22_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_22_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_22_591 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_22_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_22_661 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_22_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_22_731 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_22_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_22_801 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_22_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_22_871 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_22_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_22_941 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_22_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_23_1046 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_23_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_23_1116 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_23_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_23_1186 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_23_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_23_1256 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_23_1262 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_23_1326 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_23_1332 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_23_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_23_1396 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_23_1402 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_23_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_23_1466 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_23_1472 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_23_1536 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_23_1542 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_23_1606 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_23_1612 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_23_1676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_23_1682 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_23_1746 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_23_1752 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_23_1816 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_23_1822 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_23_1886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_23_1892 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_23_1956 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_23_1962 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_23_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_23_2026 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_23_2032 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_23_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_23_2096 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_23_2102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_23_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_23_2166 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_23_2172 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_23_2236 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_23_2242 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_23_2306 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_23_2312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_23_2376 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_23_2382 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_23_2446 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_23_2452 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_23_2516 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_23_2522 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_23_2586 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_23_2592 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_23_2624 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_23_2640 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_23_2648 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_23_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_23_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_23_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_23_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_23_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_23_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_23_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_23_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_23_556 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_23_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_23_626 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_23_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_23_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_23_696 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_23_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_23_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_23_766 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_23_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_23_836 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_23_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_23_906 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_23_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_23_976 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_23_982 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_24_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_24_1011 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_24_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_24_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_24_1081 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_24_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_24_1151 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_24_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_24_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_24_1227 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_24_1291 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_24_1297 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_24_1361 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_24_1367 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_24_1431 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_24_1437 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_24_1501 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_24_1507 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_24_1571 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_24_1577 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_24_1641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_24_1647 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_24_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_24_1711 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_24_1717 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_24_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_24_1781 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_24_1787 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_24_1851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_24_1857 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_24_1921 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_24_1927 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_24_1991 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_24_1997 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_24_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_24_2061 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_24_2067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_24_2131 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_24_2137 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_24_2201 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_24_2207 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_24_2271 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_24_2277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_24_2341 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_24_2347 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_24_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_24_2411 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_24_2417 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_24_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_24_2481 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_24_2487 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_24_2551 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_24_2557 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_24_2621 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_24_2627 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_24_2643 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_24_2651 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_24_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_24_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_24_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_24_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_24_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_24_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_24_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_24_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_24_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_24_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_24_591 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_24_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_24_661 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_24_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_24_731 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_24_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_24_801 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_24_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_24_871 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_24_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_24_941 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_24_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_25_1046 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_25_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_25_1116 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_25_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_25_1186 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_25_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_25_1256 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_25_1262 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_25_1326 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_25_1332 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_25_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_25_1396 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_25_1402 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_25_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_25_1466 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_25_1472 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_25_1536 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_25_1542 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_25_1606 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_25_1612 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_25_1676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_25_1682 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_25_1746 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_25_1752 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_25_1816 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_25_1822 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_25_1886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_25_1892 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_25_1956 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_25_1962 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_25_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_25_2026 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_25_2032 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_25_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_25_2096 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_25_2102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_25_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_25_2166 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_25_2172 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_25_2236 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_25_2242 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_25_2306 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_25_2312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_25_2376 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_25_2382 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_25_2446 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_25_2452 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_25_2516 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_25_2522 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_25_2586 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_25_2592 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_25_2624 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_25_2640 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_25_2648 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_25_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_25_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_25_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_25_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_25_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_25_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_25_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_25_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_25_556 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_25_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_25_626 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_25_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_25_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_25_696 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_25_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_25_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_25_766 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_25_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_25_836 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_25_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_25_906 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_25_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_25_976 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_25_982 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_26_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_26_1011 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_26_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_26_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_26_1081 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_26_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_26_1151 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_26_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_26_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_26_1227 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_26_1291 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_26_1297 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_26_1361 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_26_1367 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_26_1431 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_26_1437 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_26_1501 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_26_1507 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_26_1571 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_26_1577 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_26_1641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_26_1647 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_26_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_26_1711 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_26_1717 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_26_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_26_1781 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_26_1787 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_26_1851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_26_1857 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_26_1921 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_26_1927 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_26_1991 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_26_1997 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_26_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_26_2061 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_26_2067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_26_2131 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_26_2137 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_26_2201 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_26_2207 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_26_2271 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_26_2277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_26_2341 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_26_2347 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_26_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_26_2411 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_26_2417 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_26_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_26_2481 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_26_2487 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_26_2551 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_26_2557 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_26_2621 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_26_2627 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_26_2643 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_26_2651 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_26_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_26_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_26_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_26_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_26_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_26_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_26_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_26_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_26_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_26_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_26_591 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_26_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_26_661 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_26_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_26_731 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_26_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_26_801 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_26_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_26_871 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_26_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_26_941 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_26_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_27_1046 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_27_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_27_1116 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_27_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_27_1186 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_27_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_27_1256 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_27_1262 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_27_1326 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_27_1332 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_27_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_27_1396 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_27_1402 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_27_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_27_1466 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_27_1472 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_27_1536 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_27_1542 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_27_1606 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_27_1612 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_27_1676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_27_1682 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_27_1746 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_27_1752 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_27_1816 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_27_1822 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_27_1886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_27_1892 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_27_1956 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_27_1962 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_27_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_27_2026 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_27_2032 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_27_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_27_2096 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_27_2102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_27_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_27_2166 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_27_2172 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_27_2236 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_27_2242 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_27_2306 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_27_2312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_27_2376 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_27_2382 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_27_2446 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_27_2452 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_27_2516 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_27_2522 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_27_2586 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_27_2592 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_27_2624 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_27_2640 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_27_2648 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_27_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_27_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_27_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_27_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_27_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_27_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_27_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_27_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_27_556 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_27_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_27_626 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_27_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_27_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_27_696 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_27_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_27_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_27_766 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_27_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_27_836 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_27_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_27_906 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_27_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_27_976 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_27_982 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_28_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_28_1011 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_28_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_28_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_28_1081 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_28_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_28_1151 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_28_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_28_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_28_1227 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_28_1291 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_28_1297 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_28_1361 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_28_1367 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_28_1431 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_28_1437 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_28_1501 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_28_1507 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_28_1571 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_28_1577 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_28_1641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_28_1647 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_28_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_28_1711 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_28_1717 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_28_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_28_1781 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_28_1787 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_28_1851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_28_1857 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_28_1921 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_28_1927 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_28_1991 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_28_1997 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_28_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_28_2061 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_28_2067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_28_2131 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_28_2137 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_28_2201 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_28_2207 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_28_2271 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_28_2277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_28_2341 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_28_2347 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_28_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_28_2411 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_28_2417 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_28_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_28_2481 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_28_2487 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_28_2551 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_28_2557 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_28_2621 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_28_2627 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_28_2643 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_28_2651 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_28_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_28_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_28_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_28_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_28_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_28_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_28_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_28_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_28_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_28_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_28_591 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_28_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_28_661 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_28_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_28_731 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_28_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_28_801 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_28_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_28_871 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_28_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_28_941 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_28_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_29_1046 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_29_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_29_1116 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_29_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_29_1186 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_29_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_29_1256 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_29_1262 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_29_1326 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_29_1332 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_29_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_29_1396 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_29_1402 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_29_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_29_1466 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_29_1472 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_29_1536 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_29_1542 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_29_1606 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_29_1612 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_29_1676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_29_1682 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_29_1746 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_29_1752 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_29_1816 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_29_1822 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_29_1886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_29_1892 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_29_1956 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_29_1962 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_29_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_29_2026 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_29_2032 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_29_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_29_2096 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_29_2102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_29_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_29_2166 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_29_2172 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_29_2236 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_29_2242 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_29_2306 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_29_2312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_29_2376 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_29_2382 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_29_2446 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_29_2452 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_29_2516 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_29_2522 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_29_2586 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_29_2592 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_29_2624 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_29_2640 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_29_2648 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_29_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_29_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_29_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_29_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_29_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_29_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_29_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_29_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_29_556 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_29_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_29_626 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_29_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_29_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_29_696 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_29_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_29_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_29_766 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_29_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_29_836 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_29_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_29_906 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_29_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_29_976 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_29_982 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_2_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_2_1011 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_2_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_2_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_2_1081 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_2_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_2_1151 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_2_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_2_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_2_1227 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_2_1291 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_2_1297 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_2_1361 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_2_1367 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_2_1431 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_2_1437 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_2_1501 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_2_1507 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_2_1571 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_2_1577 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_2_1609 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_2_1656 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_2_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_2_1727 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_2_1731 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_2_1735 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_2_1737 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_2_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_2_1787 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_2_1821 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_2_1823 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_2_1842 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_2_1846 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_2_1874 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_2_1876 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_2_1890 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_2_1898 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_2_1921 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_2_1946 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_2_1948 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_2_1971 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_2_1991 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_2_1997 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_2_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_2_2061 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_2_2067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_2_2131 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_2_2137 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_2_2201 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_2_2207 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_2_2271 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_2_2277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_2_2341 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_2_2347 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_2_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_2_2411 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_2_2417 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_2_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_2_2481 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_2_2487 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_2_2551 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_2_2557 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_2_2621 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_2_2627 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_2_2643 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_2_2651 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_2_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_2_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_2_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_2_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_2_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_2_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_2_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_2_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_2_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_2_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_2_591 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_2_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_2_661 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_2_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_2_731 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_2_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_2_801 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_2_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_2_825 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_2_857 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_2_873 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_2_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_2_941 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_2_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_30_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_30_1011 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_30_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_30_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_30_1081 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_30_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_30_1151 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_30_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_30_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_30_1227 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_30_1291 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_30_1297 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_30_1361 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_30_1367 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_30_1431 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_30_1437 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_30_1501 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_30_1507 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_30_1571 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_30_1577 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_30_1641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_30_1647 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_30_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_30_1711 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_30_1717 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_30_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_30_1781 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_30_1787 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_30_1851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_30_1857 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_30_1921 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_30_1927 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_30_1991 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_30_1997 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_30_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_30_2061 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_30_2067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_30_2131 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_30_2137 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_30_2201 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_30_2207 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_30_2271 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_30_2277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_30_2341 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_30_2347 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_30_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_30_2411 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_30_2417 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_30_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_30_2481 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_30_2487 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_30_2551 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_30_2557 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_30_2621 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_30_2627 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_30_2643 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_30_2651 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_30_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_30_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_30_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_30_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_30_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_30_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_30_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_30_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_30_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_30_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_30_591 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_30_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_30_661 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_30_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_30_731 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_30_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_30_801 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_30_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_30_871 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_30_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_30_941 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_30_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_31_1046 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_31_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_31_1116 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_31_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_31_1186 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_31_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_31_1256 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_31_1262 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_31_1326 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_31_1332 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_31_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_31_1396 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_31_1402 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_31_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_31_1466 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_31_1472 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_31_1536 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_31_1542 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_31_1606 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_31_1612 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_31_1676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_31_1682 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_31_1746 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_31_1752 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_31_1816 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_31_1822 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_31_1886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_31_1892 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_31_1956 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_31_1962 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_31_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_31_2026 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_31_2032 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_31_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_31_2096 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_31_2102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_31_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_31_2166 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_31_2172 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_31_2236 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_31_2242 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_31_2306 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_31_2312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_31_2376 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_31_2382 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_31_2446 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_31_2452 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_31_2516 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_31_2522 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_31_2586 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_31_2592 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_31_2624 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_31_2640 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_31_2648 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_31_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_31_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_31_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_31_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_31_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_31_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_31_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_31_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_31_556 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_31_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_31_626 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_31_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_31_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_31_696 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_31_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_31_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_31_766 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_31_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_31_836 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_31_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_31_906 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_31_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_31_976 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_31_982 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_32_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_32_1011 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_32_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_32_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_32_1081 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_32_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_32_1151 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_32_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_32_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_32_1227 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_32_1291 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_32_1297 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_32_1361 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_32_1367 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_32_1431 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_32_1437 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_32_1501 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_32_1507 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_32_1571 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_32_1577 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_32_1641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_32_1647 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_32_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_32_1711 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_32_1717 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_32_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_32_1781 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_32_1787 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_32_1851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_32_1857 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_32_1921 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_32_1927 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_32_1991 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_32_1997 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_32_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_32_2061 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_32_2067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_32_2131 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_32_2137 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_32_2201 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_32_2207 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_32_2271 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_32_2277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_32_2341 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_32_2347 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_32_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_32_2411 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_32_2417 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_32_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_32_2481 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_32_2487 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_32_2551 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_32_2557 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_32_2621 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_32_2627 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_32_2643 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_32_2651 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_32_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_32_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_32_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_32_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_32_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_32_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_32_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_32_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_32_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_32_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_32_591 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_32_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_32_661 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_32_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_32_731 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_32_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_32_801 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_32_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_32_871 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_32_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_32_941 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_32_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_33_1046 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_33_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_33_1116 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_33_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_33_1186 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_33_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_33_1256 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_33_1262 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_33_1326 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_33_1332 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_33_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_33_1396 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_33_1402 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_33_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_33_1466 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_33_1472 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_33_1536 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_33_1542 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_33_1606 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_33_1612 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_33_1676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_33_1682 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_33_1746 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_33_1752 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_33_1816 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_33_1822 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_33_1886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_33_1892 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_33_1956 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_33_1962 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_33_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_33_2026 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_33_2032 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_33_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_33_2096 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_33_2102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_33_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_33_2166 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_33_2172 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_33_2236 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_33_2242 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_33_2306 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_33_2312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_33_2376 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_33_2382 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_33_2446 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_33_2452 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_33_2516 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_33_2522 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_33_2586 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_33_2592 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_33_2624 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_33_2640 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_33_2648 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_33_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_33_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_33_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_33_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_33_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_33_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_33_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_33_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_33_556 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_33_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_33_626 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_33_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_33_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_33_696 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_33_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_33_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_33_766 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_33_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_33_836 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_33_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_33_906 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_33_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_33_976 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_33_982 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_34_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_34_1011 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_34_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_34_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_34_1081 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_34_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_34_1151 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_34_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_34_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_34_1227 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_34_1291 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_34_1297 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_34_1361 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_34_1367 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_34_1431 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_34_1437 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_34_1501 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_34_1507 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_34_1571 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_34_1577 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_34_1641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_34_1647 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_34_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_34_1711 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_34_1717 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_34_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_34_1781 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_34_1787 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_34_1851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_34_1857 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_34_1921 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_34_1927 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_34_1991 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_34_1997 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_34_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_34_2061 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_34_2067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_34_2131 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_34_2137 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_34_2201 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_34_2207 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_34_2271 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_34_2277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_34_2341 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_34_2347 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_34_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_34_2411 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_34_2417 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_34_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_34_2481 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_34_2487 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_34_2551 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_34_2557 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_34_2621 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_34_2627 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_34_2643 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_34_2651 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_34_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_34_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_34_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_34_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_34_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_34_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_34_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_34_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_34_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_34_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_34_591 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_34_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_34_661 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_34_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_34_731 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_34_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_34_801 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_34_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_34_871 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_34_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_34_941 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_34_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_35_1046 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_35_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_35_1116 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_35_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_35_1186 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_35_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_35_1256 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_35_1262 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_35_1326 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_35_1332 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_35_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_35_1396 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_35_1402 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_35_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_35_1466 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_35_1472 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_35_1536 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_35_1542 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_35_1606 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_35_1612 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_35_1676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_35_1682 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_35_1746 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_35_1752 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_35_1816 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_35_1822 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_35_1886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_35_1892 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_35_1956 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_35_1962 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_35_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_35_2026 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_35_2032 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_35_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_35_2096 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_35_2102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_35_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_35_2166 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_35_2172 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_35_2236 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_35_2242 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_35_2306 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_35_2312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_35_2376 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_35_2382 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_35_2446 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_35_2452 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_35_2516 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_35_2522 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_35_2586 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_35_2592 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_35_2624 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_35_2640 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_35_2648 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_35_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_35_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_35_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_35_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_35_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_35_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_35_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_35_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_35_556 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_35_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_35_626 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_35_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_35_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_35_696 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_35_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_35_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_35_766 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_35_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_35_836 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_35_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_35_906 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_35_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_35_976 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_35_982 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_36_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_36_1011 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_36_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_36_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_36_1081 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_36_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_36_1151 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_36_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_36_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_36_1227 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_36_1291 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_36_1297 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_36_1361 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_36_1367 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_36_1431 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_36_1437 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_36_1501 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_36_1507 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_36_1571 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_36_1577 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_36_1641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_36_1647 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_36_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_36_1711 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_36_1717 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_36_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_36_1781 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_36_1787 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_36_1851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_36_1857 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_36_1921 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_36_1927 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_36_1991 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_36_1997 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_36_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_36_2061 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_36_2067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_36_2131 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_36_2137 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_36_2201 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_36_2207 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_36_2271 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_36_2277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_36_2341 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_36_2347 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_36_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_36_2411 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_36_2417 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_36_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_36_2481 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_36_2487 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_36_2551 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_36_2557 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_36_2621 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_36_2627 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_36_2643 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_36_2651 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_36_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_36_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_36_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_36_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_36_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_36_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_36_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_36_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_36_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_36_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_36_591 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_36_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_36_661 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_36_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_36_731 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_36_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_36_801 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_36_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_36_871 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_36_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_36_941 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_36_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_37_1046 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_37_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_37_1116 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_37_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_37_1186 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_37_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_37_1256 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_37_1262 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_37_1326 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_37_1332 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_37_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_37_1396 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_37_1402 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_37_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_37_1466 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_37_1472 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_37_1536 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_37_1542 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_37_1606 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_37_1612 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_37_1676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_37_1682 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_37_1746 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_37_1752 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_37_1816 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_37_1822 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_37_1886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_37_1892 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_37_1956 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_37_1962 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_37_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_37_2026 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_37_2032 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_37_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_37_2096 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_37_2102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_37_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_37_2166 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_37_2172 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_37_2236 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_37_2242 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_37_2306 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_37_2312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_37_2376 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_37_2382 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_37_2446 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_37_2452 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_37_2516 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_37_2522 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_37_2586 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_37_2592 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_37_2624 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_37_2640 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_37_2648 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_37_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_37_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_37_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_37_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_37_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_37_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_37_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_37_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_37_556 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_37_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_37_626 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_37_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_37_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_37_696 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_37_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_37_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_37_766 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_37_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_37_836 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_37_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_37_906 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_37_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_37_976 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_37_982 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_38_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_38_1011 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_38_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_38_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_38_1081 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_38_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_38_1151 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_38_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_38_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_38_1227 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_38_1291 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_38_1297 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_38_1361 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_38_1367 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_38_1431 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_38_1437 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_38_1501 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_38_1507 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_38_1571 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_38_1577 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_38_1641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_38_1647 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_38_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_38_1711 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_38_1717 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_38_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_38_1781 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_38_1787 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_38_1851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_38_1857 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_38_1921 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_38_1927 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_38_1991 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_38_1997 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_38_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_38_2061 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_38_2067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_38_2131 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_38_2137 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_38_2201 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_38_2207 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_38_2271 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_38_2277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_38_2341 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_38_2347 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_38_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_38_2411 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_38_2417 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_38_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_38_2481 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_38_2487 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_38_2551 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_38_2557 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_38_2621 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_38_2627 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_38_2643 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_38_2651 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_38_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_38_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_38_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_38_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_38_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_38_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_38_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_38_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_38_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_38_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_38_591 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_38_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_38_661 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_38_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_38_731 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_38_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_38_801 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_38_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_38_871 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_38_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_38_941 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_38_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_39_1046 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_39_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_39_1116 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_39_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_39_1186 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_39_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_39_1256 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_39_1262 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_39_1326 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_39_1332 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_39_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_39_1396 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_39_1402 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_39_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_39_1466 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_39_1472 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_39_1536 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_39_1542 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_39_1606 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_39_1612 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_39_1676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_39_1682 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_39_1746 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_39_1752 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_39_1816 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_39_1822 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_39_1886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_39_1892 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_39_1956 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_39_1962 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_39_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_39_2026 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_39_2032 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_39_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_39_2096 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_39_2102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_39_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_39_2166 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_39_2172 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_39_2236 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_39_2242 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_39_2306 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_39_2312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_39_2376 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_39_2382 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_39_2446 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_39_2452 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_39_2516 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_39_2522 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_39_2586 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_39_2592 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_39_2624 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_39_2640 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_39_2648 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_39_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_39_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_39_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_39_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_39_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_39_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_39_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_39_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_39_556 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_39_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_39_626 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_39_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_39_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_39_696 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_39_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_39_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_39_766 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_39_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_39_836 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_39_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_39_906 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_39_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_39_976 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_39_982 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_3_1046 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_3_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_3_1116 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_3_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_3_1186 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_3_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_3_1256 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_3_1262 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_3_1326 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_3_1332 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_3_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_3_1396 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_3_1402 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_3_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_3_1466 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_3_1472 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_3_1536 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_3_1542 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_3_1606 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_3_1612 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_3_1620 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_3_1664 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_3_1668 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_3_1696 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_3_1702 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_3_1736 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_3_1747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_3_1749 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_3_1807 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_3_1811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_3_1839 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_3_1843 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_3_1847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_3_1851 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_3_1855 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_3_1857 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_3_1879 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_3_1887 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_3_1889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_3_1892 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_3_1900 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_3_1902 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_3_1909 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_3_1913 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_3_1924 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_3_1928 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_3_1944 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_3_1946 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_3_1949 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_3_1957 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_3_1959 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_3_1962 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_3_1978 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_3_1982 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_3_1985 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_3_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_3_2017 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_3_2025 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_3_2029 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_3_2032 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_3_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_3_2096 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_3_2102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_3_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_3_2166 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_3_2172 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_3_2236 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_3_2242 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_3_2306 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_3_2312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_3_2376 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_3_2382 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_3_2446 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_3_2452 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_3_2516 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_3_2522 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_3_2586 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_3_2592 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_3_2624 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_3_2640 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_3_2648 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_3_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_3_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_3_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_3_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_3_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_3_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_3_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_3_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_3_556 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_3_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_3_626 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_3_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_3_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_3_696 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_3_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_3_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_3_766 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_3_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_3_836 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_3_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_3_906 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_3_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_3_976 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_3_982 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_40_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_40_1011 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_40_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_40_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_40_1081 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_40_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_40_1151 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_40_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_40_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_40_1227 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_40_1291 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_40_1297 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_40_1361 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_40_1367 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_40_1431 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_40_1437 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_40_1501 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_40_1507 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_40_1571 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_40_1577 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_40_1641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_40_1647 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_40_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_40_1711 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_40_1717 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_40_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_40_1781 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_40_1787 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_40_1851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_40_1857 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_40_1921 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_40_1927 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_40_1991 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_40_1997 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_40_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_40_2061 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_40_2067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_40_2131 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_40_2137 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_40_2201 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_40_2207 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_40_2271 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_40_2277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_40_2341 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_40_2347 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_40_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_40_2411 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_40_2417 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_40_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_40_2481 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_40_2487 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_40_2551 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_40_2557 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_40_2621 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_40_2627 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_40_2643 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_40_2651 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_40_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_40_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_40_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_40_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_40_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_40_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_40_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_40_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_40_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_40_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_40_591 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_40_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_40_661 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_40_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_40_731 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_40_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_40_801 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_40_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_40_871 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_40_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_40_941 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_40_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_41_1046 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_41_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_41_1116 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_41_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_41_1186 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_41_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_41_1256 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_41_1262 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_41_1326 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_41_1332 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_41_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_41_1396 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_41_1402 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_41_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_41_1466 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_41_1472 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_41_1536 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_41_1542 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_41_1606 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_41_1612 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_41_1676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_41_1682 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_41_1746 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_41_1752 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_41_1816 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_41_1822 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_41_1886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_41_1892 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_41_1956 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_41_1962 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_41_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_41_2026 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_41_2032 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_41_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_41_2096 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_41_2102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_41_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_41_2166 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_41_2172 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_41_2236 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_41_2242 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_41_2306 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_41_2312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_41_2376 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_41_2382 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_41_2446 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_41_2452 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_41_2516 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_41_2522 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_41_2586 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_41_2592 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_41_2624 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_41_2640 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_41_2648 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_41_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_41_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_41_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_41_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_41_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_41_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_41_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_41_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_41_556 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_41_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_41_626 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_41_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_41_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_41_696 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_41_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_41_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_41_766 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_41_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_41_836 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_41_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_41_906 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_41_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_41_976 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_41_982 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_42_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_42_1011 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_42_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_42_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_42_1081 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_42_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_42_1151 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_42_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_42_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_42_1227 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_42_1291 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_42_1297 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_42_1361 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_42_1367 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_42_1431 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_42_1437 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_42_1501 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_42_1507 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_42_1571 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_42_1577 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_42_1641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_42_1647 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_42_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_42_1711 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_42_1717 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_42_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_42_1781 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_42_1787 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_42_1851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_42_1857 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_42_1921 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_42_1927 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_42_1991 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_42_1997 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_42_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_42_2061 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_42_2067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_42_2131 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_42_2137 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_42_2201 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_42_2207 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_42_2271 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_42_2277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_42_2341 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_42_2347 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_42_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_42_2411 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_42_2417 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_42_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_42_2481 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_42_2487 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_42_2551 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_42_2557 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_42_2621 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_42_2627 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_42_2643 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_42_2651 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_42_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_42_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_42_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_42_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_42_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_42_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_42_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_42_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_42_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_42_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_42_591 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_42_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_42_661 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_42_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_42_731 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_42_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_42_801 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_42_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_42_871 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_42_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_42_941 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_42_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_43_1046 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_43_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_43_1116 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_43_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_43_1186 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_43_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_43_1256 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_43_1262 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_43_1326 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_43_1332 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_43_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_43_1396 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_43_1402 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_43_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_43_1466 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_43_1472 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_43_1536 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_43_1542 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_43_1606 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_43_1612 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_43_1676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_43_1682 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_43_1746 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_43_1752 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_43_1816 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_43_1822 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_43_1886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_43_1892 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_43_1956 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_43_1962 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_43_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_43_2026 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_43_2032 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_43_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_43_2096 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_43_2102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_43_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_43_2166 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_43_2172 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_43_2236 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_43_2242 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_43_2306 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_43_2312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_43_2376 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_43_2382 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_43_2446 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_43_2452 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_43_2516 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_43_2522 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_43_2586 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_43_2592 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_43_2624 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_43_2640 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_43_2648 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_43_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_43_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_43_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_43_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_43_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_43_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_43_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_43_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_43_556 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_43_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_43_626 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_43_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_43_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_43_696 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_43_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_43_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_43_766 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_43_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_43_836 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_43_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_43_906 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_43_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_43_976 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_43_982 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_44_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_44_1011 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_44_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_44_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_44_1081 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_44_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_44_1151 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_44_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_44_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_44_1227 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_44_1291 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_44_1297 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_44_1361 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_44_1367 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_44_1431 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_44_1437 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_44_1501 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_44_1507 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_44_1571 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_44_1577 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_44_1641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_44_1647 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_44_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_44_1711 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_44_1717 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_44_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_44_1781 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_44_1787 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_44_1851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_44_1857 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_44_1921 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_44_1927 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_44_1991 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_44_1997 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_44_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_44_2061 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_44_2067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_44_2131 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_44_2137 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_44_2201 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_44_2207 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_44_2271 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_44_2277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_44_2341 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_44_2347 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_44_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_44_2411 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_44_2417 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_44_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_44_2481 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_44_2487 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_44_2551 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_44_2557 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_44_2621 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_44_2627 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_44_2643 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_44_2651 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_44_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_44_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_44_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_44_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_44_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_44_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_44_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_44_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_44_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_44_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_44_591 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_44_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_44_661 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_44_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_44_731 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_44_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_44_801 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_44_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_44_871 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_44_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_44_941 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_44_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_45_1046 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_45_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_45_1116 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_45_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_45_1186 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_45_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_45_1256 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_45_1262 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_45_1326 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_45_1332 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_45_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_45_1396 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_45_1402 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_45_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_45_1466 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_45_1472 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_45_1536 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_45_1542 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_45_1606 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_45_1612 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_45_1676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_45_1682 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_45_1746 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_45_1752 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_45_1816 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_45_1822 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_45_1886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_45_1892 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_45_1956 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_45_1962 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_45_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_45_2026 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_45_2032 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_45_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_45_2096 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_45_2102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_45_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_45_2166 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_45_2172 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_45_2236 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_45_2242 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_45_2306 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_45_2312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_45_2376 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_45_2382 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_45_2446 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_45_2452 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_45_2516 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_45_2522 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_45_2586 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_45_2592 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_45_2624 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_45_2640 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_45_2648 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_45_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_45_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_45_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_45_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_45_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_45_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_45_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_45_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_45_556 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_45_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_45_626 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_45_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_45_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_45_696 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_45_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_45_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_45_766 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_45_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_45_836 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_45_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_45_906 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_45_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_45_976 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_45_982 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_46_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_46_1011 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_46_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_46_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_46_1081 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_46_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_46_1151 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_46_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_46_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_46_1227 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_46_1291 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_46_1297 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_46_1361 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_46_1367 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_46_1431 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_46_1437 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_46_1501 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_46_1507 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_46_1571 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_46_1577 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_46_1641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_46_1647 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_46_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_46_1711 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_46_1717 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_46_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_46_1781 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_46_1787 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_46_1851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_46_1857 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_46_1921 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_46_1927 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_46_1991 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_46_1997 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_46_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_46_2061 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_46_2067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_46_2131 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_46_2137 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_46_2201 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_46_2207 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_46_2271 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_46_2277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_46_2341 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_46_2347 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_46_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_46_2411 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_46_2417 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_46_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_46_2481 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_46_2487 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_46_2551 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_46_2557 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_46_2621 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_46_2627 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_46_2643 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_46_2651 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_46_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_46_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_46_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_46_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_46_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_46_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_46_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_46_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_46_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_46_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_46_591 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_46_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_46_661 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_46_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_46_731 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_46_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_46_801 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_46_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_46_871 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_46_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_46_941 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_46_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_47_1046 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_47_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_47_1116 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_47_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_47_1186 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_47_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_47_1256 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_47_1262 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_47_1326 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_47_1332 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_47_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_47_1396 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_47_1402 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_47_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_47_1466 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_47_1472 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_47_1536 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_47_1542 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_47_1606 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_47_1612 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_47_1676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_47_1682 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_47_1746 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_47_1752 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_47_1816 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_47_1822 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_47_1886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_47_1892 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_47_1956 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_47_1962 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_47_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_47_2026 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_47_2032 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_47_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_47_2096 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_47_2102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_47_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_47_2166 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_47_2172 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_47_2236 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_47_2242 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_47_2306 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_47_2312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_47_2376 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_47_2382 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_47_2446 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_47_2452 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_47_2516 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_47_2522 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_47_2586 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_47_2592 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_47_2624 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_47_2640 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_47_2648 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_47_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_47_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_47_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_47_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_47_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_47_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_47_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_47_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_47_556 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_47_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_47_626 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_47_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_47_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_47_696 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_47_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_47_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_47_766 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_47_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_47_836 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_47_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_47_906 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_47_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_47_976 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_47_982 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_48_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_48_1011 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_48_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_48_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_48_1081 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_48_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_48_1151 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_48_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_48_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_48_1227 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_48_1291 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_48_1297 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_48_1361 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_48_1367 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_48_1431 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_48_1437 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_48_1501 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_48_1507 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_48_1571 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_48_1577 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_48_1641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_48_1647 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_48_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_48_1711 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_48_1717 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_48_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_48_1781 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_48_1787 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_48_1851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_48_1857 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_48_1921 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_48_1927 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_48_1991 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_48_1997 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_48_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_48_2061 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_48_2067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_48_2131 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_48_2137 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_48_2201 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_48_2207 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_48_2271 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_48_2277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_48_2341 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_48_2347 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_48_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_48_2411 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_48_2417 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_48_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_48_2481 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_48_2487 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_48_2551 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_48_2557 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_48_2621 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_48_2627 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_48_2643 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_48_2651 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_48_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_48_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_48_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_48_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_48_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_48_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_48_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_48_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_48_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_48_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_48_591 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_48_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_48_661 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_48_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_48_731 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_48_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_48_801 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_48_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_48_871 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_48_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_48_941 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_48_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_49_1046 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_49_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_49_1116 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_49_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_49_1186 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_49_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_49_1256 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_49_1262 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_49_1326 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_49_1332 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_49_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_49_1396 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_49_1402 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_49_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_49_1466 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_49_1472 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_49_1536 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_49_1542 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_49_1606 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_49_1612 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_49_1676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_49_1682 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_49_1746 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_49_1752 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_49_1816 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_49_1822 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_49_1886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_49_1892 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_49_1956 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_49_1962 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_49_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_49_2026 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_49_2032 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_49_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_49_2096 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_49_2102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_49_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_49_2166 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_49_2172 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_49_2236 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_49_2242 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_49_2306 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_49_2312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_49_2376 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_49_2382 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_49_2446 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_49_2452 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_49_2516 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_49_2522 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_49_2586 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_49_2592 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_49_2624 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_49_2640 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_49_2648 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_49_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_49_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_49_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_49_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_49_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_49_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_49_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_49_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_49_556 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_49_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_49_626 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_49_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_49_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_49_696 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_49_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_49_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_49_766 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_49_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_49_836 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_49_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_49_906 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_49_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_49_976 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_49_982 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_4_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_4_1011 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_4_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_4_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_4_1081 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_4_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_4_1151 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_4_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_4_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_4_1227 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_4_1291 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_4_1297 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_4_1361 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_4_1367 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_4_1431 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_4_1437 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_4_1501 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_4_1507 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_4_1571 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_4_1577 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_4_1609 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_4_1625 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_4_1629 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_4_1637 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_4_1647 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_4_1651 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_4_1653 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_4_1656 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_4_1707 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_4_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_4_1711 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_4_1717 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_4_1721 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_4_1725 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_4_1733 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_4_1735 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_4_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_4_1834 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_4_1838 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_4_1842 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_4_1846 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_4_1854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_4_1857 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_4_1889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_4_1893 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_4_1900 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_4_1916 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_4_1924 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_4_1941 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_4_1945 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_4_1977 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_4_1993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_4_1997 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_4_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_4_2061 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_4_2067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_4_2131 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_4_2137 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_4_2201 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_4_2207 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_4_2271 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_4_2277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_4_2341 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_4_2347 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_4_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_4_2411 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_4_2417 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_4_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_4_2481 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_4_2487 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_4_2551 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_4_2557 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_4_2621 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_4_2627 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_4_2643 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_4_2651 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_4_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_4_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_4_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_4_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_4_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_4_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_4_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_4_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_4_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_4_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_4_591 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_4_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_4_661 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_4_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_4_731 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_4_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_4_801 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_4_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_4_871 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_4_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_4_941 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_4_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_50_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_50_1011 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_50_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_50_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_50_1081 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_50_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_50_1151 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_50_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_50_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_50_1227 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_50_1291 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_50_1297 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_50_1361 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_50_1367 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_50_1431 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_50_1437 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_50_1501 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_50_1507 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_50_1571 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_50_1577 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_50_1641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_50_1647 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_50_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_50_1711 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_50_1717 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_50_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_50_1781 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_50_1787 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_50_1851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_50_1857 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_50_1921 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_50_1927 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_50_1991 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_50_1997 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_50_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_50_2061 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_50_2067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_50_2131 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_50_2137 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_50_2201 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_50_2207 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_50_2271 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_50_2277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_50_2341 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_50_2347 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_50_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_50_2411 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_50_2417 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_50_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_50_2481 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_50_2487 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_50_2551 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_50_2557 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_50_2621 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_50_2627 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_50_2643 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_50_2651 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_50_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_50_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_50_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_50_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_50_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_50_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_50_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_50_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_50_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_50_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_50_591 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_50_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_50_661 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_50_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_50_731 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_50_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_50_801 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_50_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_50_871 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_50_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_50_941 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_50_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_51_1046 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_51_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_51_1116 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_51_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_51_1186 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_51_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_51_1256 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_51_1262 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_51_1326 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_51_1332 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_51_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_51_1396 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_51_1402 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_51_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_51_1466 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_51_1472 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_51_1536 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_51_1542 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_51_1606 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_51_1612 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_51_1676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_51_1682 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_51_1746 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_51_1752 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_51_1816 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_51_1822 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_51_1886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_51_1892 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_51_1956 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_51_1962 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_51_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_51_2026 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_51_2032 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_51_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_51_2096 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_51_2102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_51_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_51_2166 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_51_2172 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_51_2236 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_51_2242 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_51_2306 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_51_2312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_51_2376 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_51_2382 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_51_2446 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_51_2452 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_51_2516 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_51_2522 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_51_2586 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_51_2592 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_51_2624 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_51_2640 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_51_2648 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_51_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_51_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_51_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_51_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_51_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_51_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_51_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_51_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_51_556 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_51_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_51_626 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_51_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_51_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_51_696 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_51_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_51_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_51_766 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_51_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_51_836 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_51_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_51_906 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_51_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_51_976 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_51_982 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_52_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_52_1011 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_52_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_52_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_52_1081 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_52_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_52_1151 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_52_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_52_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_52_1227 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_52_1291 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_52_1297 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_52_1361 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_52_1367 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_52_1431 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_52_1437 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_52_1501 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_52_1507 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_52_1571 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_52_1577 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_52_1641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_52_1647 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_52_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_52_1711 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_52_1717 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_52_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_52_1781 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_52_1787 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_52_1851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_52_1857 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_52_1921 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_52_1927 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_52_1991 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_52_1997 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_52_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_52_2061 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_52_2067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_52_2131 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_52_2137 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_52_2201 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_52_2207 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_52_2271 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_52_2277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_52_2341 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_52_2347 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_52_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_52_2411 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_52_2417 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_52_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_52_2481 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_52_2487 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_52_2551 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_52_2557 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_52_2621 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_52_2627 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_52_2643 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_52_2651 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_52_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_52_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_52_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_52_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_52_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_52_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_52_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_52_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_52_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_52_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_52_591 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_52_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_52_661 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_52_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_52_731 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_52_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_52_801 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_52_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_52_871 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_52_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_52_941 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_52_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_53_1046 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_53_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_53_1116 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_53_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_53_1186 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_53_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_53_1256 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_53_1262 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_53_1326 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_53_1332 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_53_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_53_1396 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_53_1402 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_53_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_53_1466 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_53_1472 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_53_1536 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_53_1542 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_53_1606 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_53_1612 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_53_1676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_53_1682 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_53_1746 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_53_1752 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_53_1816 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_53_1822 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_53_1886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_53_1892 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_53_1956 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_53_1962 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_53_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_53_2026 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_53_2032 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_53_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_53_2096 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_53_2102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_53_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_53_2166 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_53_2172 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_53_2236 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_53_2242 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_53_2306 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_53_2312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_53_2376 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_53_2382 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_53_2446 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_53_2452 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_53_2516 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_53_2522 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_53_2586 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_53_2592 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_53_2624 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_53_2640 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_53_2648 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_53_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_53_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_53_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_53_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_53_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_53_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_53_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_53_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_53_556 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_53_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_53_626 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_53_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_53_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_53_696 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_53_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_53_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_53_766 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_53_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_53_836 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_53_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_53_906 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_53_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_53_976 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_53_982 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_54_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_54_1011 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_54_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_54_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_54_1081 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_54_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_54_1151 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_54_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_54_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_54_1227 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_54_1291 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_54_1297 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_54_1361 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_54_1367 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_54_1431 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_54_1437 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_54_1501 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_54_1507 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_54_1571 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_54_1577 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_54_1641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_54_1647 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_54_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_54_1711 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_54_1717 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_54_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_54_1781 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_54_1787 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_54_1851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_54_1857 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_54_1921 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_54_1927 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_54_1991 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_54_1997 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_54_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_54_2061 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_54_2067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_54_2131 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_54_2137 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_54_2201 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_54_2207 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_54_2271 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_54_2277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_54_2341 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_54_2347 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_54_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_54_2411 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_54_2417 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_54_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_54_2481 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_54_2487 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_54_2551 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_54_2557 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_54_2621 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_54_2627 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_54_2643 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_54_2651 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_54_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_54_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_54_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_54_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_54_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_54_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_54_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_54_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_54_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_54_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_54_591 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_54_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_54_661 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_54_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_54_731 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_54_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_54_801 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_54_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_54_871 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_54_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_54_941 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_54_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_55_1046 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_55_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_55_1116 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_55_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_55_1186 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_55_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_55_1256 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_55_1262 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_55_1326 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_55_1332 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_55_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_55_1396 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_55_1402 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_55_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_55_1466 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_55_1472 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_55_1536 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_55_1542 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_55_1606 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_55_1612 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_55_1676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_55_1682 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_55_1746 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_55_1752 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_55_1816 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_55_1822 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_55_1886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_55_1892 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_55_1956 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_55_1962 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_55_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_55_2026 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_55_2032 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_55_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_55_2096 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_55_2102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_55_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_55_2166 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_55_2172 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_55_2236 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_55_2242 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_55_2306 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_55_2312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_55_2376 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_55_2382 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_55_2446 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_55_2452 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_55_2516 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_55_2522 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_55_2586 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_55_2592 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_55_2624 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_55_2640 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_55_2648 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_55_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_55_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_55_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_55_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_55_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_55_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_55_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_55_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_55_556 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_55_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_55_626 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_55_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_55_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_55_696 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_55_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_55_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_55_766 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_55_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_55_836 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_55_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_55_906 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_55_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_55_976 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_55_982 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_56_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_56_1011 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_56_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_56_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_56_1081 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_56_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_56_1151 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_56_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_56_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_56_1227 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_56_1291 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_56_1297 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_56_1361 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_56_1367 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_56_1431 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_56_1437 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_56_1501 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_56_1507 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_56_1571 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_56_1577 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_56_1641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_56_1647 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_56_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_56_1711 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_56_1717 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_56_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_56_1781 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_56_1787 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_56_1851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_56_1857 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_56_1921 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_56_1927 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_56_1991 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_56_1997 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_56_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_56_2061 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_56_2067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_56_2131 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_56_2137 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_56_2201 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_56_2207 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_56_2271 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_56_2277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_56_2341 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_56_2347 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_56_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_56_2411 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_56_2417 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_56_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_56_2481 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_56_2487 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_56_2551 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_56_2557 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_56_2621 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_56_2627 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_56_2643 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_56_2651 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_56_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_56_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_56_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_56_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_56_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_56_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_56_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_56_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_56_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_56_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_56_591 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_56_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_56_661 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_56_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_56_731 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_56_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_56_801 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_56_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_56_871 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_56_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_56_941 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_56_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_57_1046 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_57_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_57_1116 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_57_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_57_1186 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_57_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_57_1256 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_57_1262 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_57_1326 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_57_1332 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_57_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_57_1396 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_57_1402 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_57_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_57_1466 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_57_1472 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_57_1536 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_57_1542 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_57_1606 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_57_1612 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_57_1676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_57_1682 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_57_1746 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_57_1752 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_57_1816 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_57_1822 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_57_1886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_57_1892 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_57_1956 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_57_1962 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_57_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_57_2026 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_57_2032 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_57_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_57_2096 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_57_2102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_57_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_57_2166 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_57_2172 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_57_2236 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_57_2242 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_57_2306 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_57_2312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_57_2376 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_57_2382 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_57_2446 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_57_2452 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_57_2516 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_57_2522 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_57_2586 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_57_2592 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_57_2624 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_57_2640 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_57_2648 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_57_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_57_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_57_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_57_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_57_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_57_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_57_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_57_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_57_556 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_57_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_57_626 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_57_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_57_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_57_696 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_57_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_57_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_57_766 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_57_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_57_836 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_57_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_57_906 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_57_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_57_976 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_57_982 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_58_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_58_1011 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_58_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_58_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_58_1081 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_58_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_58_1151 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_58_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_58_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_58_1227 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_58_1291 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_58_1297 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_58_1361 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_58_1367 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_58_1431 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_58_1437 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_58_1501 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_58_1507 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_58_1571 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_58_1577 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_58_1641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_58_1647 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_58_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_58_1711 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_58_1717 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_58_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_58_1781 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_58_1787 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_58_1851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_58_1857 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_58_1921 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_58_1927 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_58_1991 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_58_1997 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_58_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_58_2061 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_58_2067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_58_2131 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_58_2137 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_58_2201 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_58_2207 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_58_2271 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_58_2277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_58_2341 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_58_2347 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_58_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_58_2411 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_58_2417 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_58_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_58_2481 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_58_2487 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_58_2551 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_58_2557 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_58_2621 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_58_2627 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_58_2643 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_58_2651 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_58_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_58_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_58_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_58_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_58_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_58_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_58_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_58_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_58_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_58_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_58_591 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_58_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_58_661 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_58_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_58_731 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_58_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_58_801 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_58_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_58_871 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_58_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_58_941 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_58_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_59_1046 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_59_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_59_1116 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_59_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_59_1186 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_59_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_59_1256 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_59_1262 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_59_1326 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_59_1332 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_59_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_59_1396 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_59_1402 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_59_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_59_1466 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_59_1472 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_59_1536 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_59_1542 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_59_1606 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_59_1612 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_59_1676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_59_1682 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_59_1746 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_59_1752 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_59_1816 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_59_1822 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_59_1886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_59_1892 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_59_1956 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_59_1962 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_59_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_59_2026 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_59_2032 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_59_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_59_2096 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_59_2102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_59_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_59_2166 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_59_2172 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_59_2236 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_59_2242 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_59_2306 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_59_2312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_59_2376 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_59_2382 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_59_2446 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_59_2452 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_59_2516 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_59_2522 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_59_2586 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_59_2592 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_59_2624 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_59_2640 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_59_2648 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_59_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_59_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_59_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_59_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_59_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_59_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_59_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_59_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_59_556 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_59_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_59_626 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_59_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_59_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_59_696 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_59_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_59_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_59_766 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_59_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_59_836 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_59_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_59_906 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_59_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_59_976 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_59_982 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_5_1046 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_5_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_5_1116 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_5_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_5_1186 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_5_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_5_1256 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_5_1262 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_5_1326 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_5_1332 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_5_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_5_1396 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_5_1402 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_5_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_5_1466 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_5_1472 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_5_1536 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_5_1542 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_5_1606 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_5_1612 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_5_1628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_5_1636 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_5_1638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_5_1692 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_5_1696 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_5_1700 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_5_1736 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_5_1740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_5_1748 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_5_1762 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_5_1764 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_5_1767 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_5_1811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_5_1813 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_5_1828 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_5_1832 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_5_1841 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_5_1857 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_5_1886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_5_1892 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_5_1896 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_5_1906 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_5_1925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_5_1957 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_5_1959 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_5_1962 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_5_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_5_2026 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_5_2032 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_5_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_5_2096 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_5_2102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_5_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_5_2166 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_5_2172 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_5_2236 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_5_2242 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_5_2306 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_5_2312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_5_2376 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_5_2382 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_5_2446 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_5_2452 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_5_2516 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_5_2522 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_5_2586 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_5_2592 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_5_2624 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_5_2640 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_5_2648 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_5_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_5_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_5_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_5_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_5_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_5_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_5_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_5_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_5_556 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_5_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_5_626 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_5_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_5_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_5_696 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_5_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_5_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_5_766 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_5_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_5_836 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_5_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_5_906 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_5_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_5_976 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_5_982 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_60_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_60_1011 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_60_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_60_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_60_1081 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_60_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_60_1151 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_60_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_60_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_60_1227 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_60_1291 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_60_1297 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_60_1361 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_60_1367 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_60_1431 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_60_1437 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_60_1501 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_60_1507 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_60_1571 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_60_1577 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_60_1641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_60_1647 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_60_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_60_1711 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_60_1717 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_60_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_60_1781 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_60_1787 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_60_1851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_60_1857 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_60_1921 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_60_1927 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_60_1991 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_60_1997 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_60_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_60_2061 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_60_2067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_60_2131 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_60_2137 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_60_2201 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_60_2207 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_60_2271 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_60_2277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_60_2341 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_60_2347 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_60_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_60_2411 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_60_2417 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_60_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_60_2481 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_60_2487 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_60_2551 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_60_2557 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_60_2621 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_60_2627 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_60_2643 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_60_2651 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_60_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_60_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_60_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_60_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_60_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_60_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_60_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_60_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_60_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_60_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_60_591 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_60_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_60_661 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_60_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_60_731 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_60_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_60_801 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_60_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_60_871 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_60_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_60_941 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_60_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_61_1046 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_61_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_61_1116 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_61_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_61_1186 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_61_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_61_1256 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_61_1262 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_61_1326 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_61_1332 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_61_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_61_1396 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_61_1402 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_61_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_61_1466 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_61_1472 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_61_1536 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_61_1542 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_61_1606 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_61_1612 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_61_1676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_61_1682 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_61_1746 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_61_1752 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_61_1816 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_61_1822 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_61_1886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_61_1892 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_61_1956 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_61_1962 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_61_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_61_2026 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_61_2032 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_61_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_61_2096 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_61_2102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_61_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_61_2166 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_61_2172 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_61_2236 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_61_2242 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_61_2306 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_61_2312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_61_2376 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_61_2382 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_61_2446 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_61_2452 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_61_2516 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_61_2522 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_61_2586 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_61_2592 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_61_2624 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_61_2640 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_61_2648 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_61_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_61_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_61_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_61_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_61_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_61_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_61_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_61_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_61_556 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_61_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_61_626 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_61_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_61_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_61_696 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_61_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_61_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_61_766 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_61_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_61_836 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_61_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_61_906 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_61_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_61_976 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_61_982 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_62_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_62_1011 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_62_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_62_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_62_1081 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_62_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_62_1151 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_62_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_62_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_62_1227 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_62_1291 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_62_1297 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_62_1361 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_62_1367 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_62_1431 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_62_1437 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_62_1501 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_62_1507 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_62_1571 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_62_1577 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_62_1641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_62_1647 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_62_1651 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_62_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_62_1717 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_62_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_62_1781 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_62_1787 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_62_1851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_62_1857 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_62_1921 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_62_1927 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_62_1991 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_62_1997 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_62_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_62_2061 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_62_2067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_62_2131 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_62_2137 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_62_2201 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_62_2207 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_62_2271 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_62_2277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_62_2341 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_62_2347 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_62_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_62_2411 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_62_2417 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_62_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_62_2481 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_62_2487 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_62_2551 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_62_2557 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_62_2621 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_62_2627 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_62_2643 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_62_2651 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_62_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_62_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_62_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_62_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_62_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_62_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_62_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_62_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_62_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_62_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_62_591 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_62_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_62_661 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_62_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_62_731 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_62_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_62_801 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_62_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_62_871 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_62_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_62_941 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_62_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_63_1046 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_63_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_63_1116 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_63_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_63_1186 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_63_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_63_1256 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_63_1262 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_63_1326 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_63_1332 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_63_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_63_1396 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_63_1402 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_63_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_63_1466 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_63_1472 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_63_1536 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_63_1542 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_63_1606 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_63_1612 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_63_1645 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_63_1649 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_63_1682 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_63_1746 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_63_1752 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_63_1816 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_63_1822 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_63_1886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_63_1892 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_63_1956 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_63_1962 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_63_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_63_2026 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_63_2032 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_63_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_63_2096 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_63_2102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_63_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_63_2166 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_63_2172 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_63_2236 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_63_2242 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_63_2306 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_63_2312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_63_2376 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_63_2382 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_63_2446 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_63_2452 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_63_2516 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_63_2522 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_63_2586 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_63_2592 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_63_2624 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_63_2640 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_63_2648 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_63_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_63_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_63_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_63_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_63_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_63_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_63_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_63_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_63_556 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_63_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_63_626 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_63_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_63_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_63_696 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_63_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_63_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_63_766 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_63_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_63_836 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_63_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_63_906 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_63_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_63_976 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_63_982 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_64_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_64_1011 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_64_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_64_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_64_1081 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_64_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_64_1119 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_64_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_64_1153 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_64_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_64_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_64_1227 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_64_1259 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_64_1275 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_64_1293 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_64_1297 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_64_1329 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_64_1343 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_64_1359 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_64_1363 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_64_1367 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_64_1431 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_64_1487 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_64_1503 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_64_1507 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_64_1571 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_64_1627 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_64_1643 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_64_1647 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_64_1663 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_64_1671 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_64_1675 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_64_1677 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_64_1680 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_64_1684 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_64_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_64_1717 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_64_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_64_1781 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_64_1787 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_64_1851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_64_1857 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_64_1921 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_64_1927 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_64_1991 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_64_1997 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_64_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_64_2061 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_64_2067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_64_2131 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_64_2137 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_64_2201 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_64_2207 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_64_2271 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_64_2277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_64_2341 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_64_2347 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_64_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_64_2411 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_64_2417 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_64_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_64_2481 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_64_2487 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_64_2551 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_64_2557 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_64_2621 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_64_2627 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_64_2643 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_64_2651 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_64_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_64_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_64_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_64_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_64_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_64_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_64_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_64_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_64_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_64_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_64_591 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_64_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_64_661 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_64_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_64_731 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_64_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_64_801 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_64_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_64_871 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_64_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_64_941 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_64_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_65_1046 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_65_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_65_1116 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_65_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_65_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_65_1142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_65_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_65_1177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_65_1185 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_65_1189 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_65_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_65_1234 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_65_1238 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_65_1249 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_65_1257 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_65_1259 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_65_1262 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_65_1278 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_65_1282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_65_1313 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_65_1317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_65_1325 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_65_1327 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_65_1332 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_65_1334 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_65_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_65_1364 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_65_1380 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_65_1382 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_65_1393 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_65_1397 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_65_1399 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_65_1402 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_65_1418 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_65_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_65_1426 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_65_1428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_65_1439 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_65_1455 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_65_1463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_65_1467 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_65_1469 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_65_1472 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_65_1476 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_65_1478 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_65_1489 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_65_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_65_1532 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_65_1542 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_65_1606 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_65_1612 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_65_1620 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_65_1652 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_65_1668 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_65_1676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_65_1682 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_65_1690 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_65_1694 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_65_1696 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_65_1728 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_65_1744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_65_1748 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_65_1752 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_65_1816 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_65_1822 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_65_1886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_65_1892 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_65_1956 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_65_1962 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_65_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_65_2026 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_65_2032 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_65_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_65_2096 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_65_2102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_65_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_65_2166 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_65_2172 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_65_2236 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_65_2242 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_65_2306 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_65_2312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_65_2376 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_65_2382 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_65_2446 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_65_2452 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_65_2516 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_65_2522 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_65_2586 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_65_2592 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_65_2624 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_65_2640 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_65_2648 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_65_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_65_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_65_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_65_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_65_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_65_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_65_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_65_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_65_556 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_65_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_65_626 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_65_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_65_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_65_696 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_65_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_65_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_65_766 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_65_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_65_836 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_65_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_65_906 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_65_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_65_976 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_65_982 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_66_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_66_1011 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_66_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_66_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_66_1081 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_66_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_66_1151 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_66_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_66_1189 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_66_1191 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_66_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_66_1227 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_66_1235 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_66_1239 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_66_1270 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_66_1274 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_66_1290 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_66_1294 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_66_1297 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_66_1301 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_66_1303 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_66_1354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_66_1358 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_66_1362 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_66_1364 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_66_1367 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_66_1414 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_66_1430 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_66_1432 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_66_1466 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_66_1474 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_66_1507 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_66_1511 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_66_1519 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_66_1523 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_66_1553 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_66_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_66_1573 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_66_1577 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_66_1585 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_66_1618 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_66_1622 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_66_1638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_66_1642 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_66_1644 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_66_1660 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_66_1664 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_66_1697 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_66_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_66_1713 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_66_1717 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_66_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_66_1781 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_66_1787 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_66_1851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_66_1857 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_66_1921 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_66_1927 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_66_1991 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_66_1997 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_66_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_66_2061 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_66_2067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_66_2131 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_66_2137 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_66_2201 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_66_2207 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_66_2271 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_66_2277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_66_2341 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_66_2347 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_66_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_66_2411 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_66_2417 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_66_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_66_2481 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_66_2487 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_66_2551 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_66_2557 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_66_2621 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_66_2627 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_66_2643 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_66_2651 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_66_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_66_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_66_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_66_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_66_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_66_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_66_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_66_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_66_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_66_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_66_591 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_66_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_66_629 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_66_657 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_66_661 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_66_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_66_731 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_66_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_66_801 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_66_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_66_871 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_66_903 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_66_907 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_66_939 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_66_943 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_66_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_67_1004 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_67_1012 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_67_1016 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_67_1030 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_67_1046 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_67_1056 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_67_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_67_1071 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_67_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_67_1090 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_67_110 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_67_1106 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_67_1108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_67_1117 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_67_1121 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_67_1124 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_67_1140 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_67_1148 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_67_1152 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_67_1158 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_67_1165 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_67_1181 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_67_1189 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_67_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_67_1200 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_67_1204 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_67_1213 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_67_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_67_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_67_1226 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_67_1242 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_67_1250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_67_1254 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_67_126 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_67_1266 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_67_1282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_67_1290 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_67_1294 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_67_1298 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_67_1300 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_67_1309 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_67_1325 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_67_1328 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_67_134 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_67_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_67_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_67_1357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_67_1359 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_67_1362 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_67_1378 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_67_138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_67_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_67_1390 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_67_1396 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_67_1398 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_67_1405 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_67_1421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_67_1425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_67_1427 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_67_1430 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_67_1438 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_67_1442 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_67_1444 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_67_1453 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_67_146 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_67_1461 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_67_1464 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_67_148 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_67_1480 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_67_1488 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_67_1492 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_67_1504 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_67_1520 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_67_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_67_1532 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_67_1540 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_67_1549 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_67_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_67_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_67_1563 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_67_1566 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_67_1582 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_67_1586 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_67_1588 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_67_1597 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_67_1600 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_67_161 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_67_1634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_67_1636 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_67_1645 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_67_1661 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_67_1663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_67_169 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_67_1702 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_67_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_67_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_67_1722 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_67_1730 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_67_1742 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_67_1758 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_67_1766 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_67_1770 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_67_1774 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_67_1804 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_67_1808 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_67_1824 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_67_1832 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_67_1864 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_67_1868 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_67_1872 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_67_1876 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_67_188 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_67_1885 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_67_1901 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_67_1903 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_67_1906 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_67_1922 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_67_1924 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_67_1933 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_67_1937 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_67_1940 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_67_1956 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_67_196 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_67_1964 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_67_1968 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_67_1974 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_67_1981 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_67_1997 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_67_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_67_200 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_67_2005 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_67_2008 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_67_2016 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_67_2020 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_67_2029 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_67_2037 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_67_2039 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_67_2042 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_67_2058 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_67_2066 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_67_2070 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_67_2082 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_67_2098 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_67_2106 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_67_2110 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_67_2114 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_67_2116 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_67_2127 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_67_2135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_67_2139 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_67_214 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_67_2141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_67_2144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_67_2160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_67_2164 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_67_2175 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_67_2178 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_67_2194 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_67_2202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_67_2206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_67_2212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_67_2214 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_67_2223 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_67_2239 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_67_2243 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_67_2246 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_67_2254 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_67_2258 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_67_2260 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_67_2277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_67_2280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_67_2296 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_67_230 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_67_2304 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_67_2308 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_67_2328 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_67_2344 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_67_2348 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_67_2356 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_67_2373 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_67_2377 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_67_2379 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_67_2382 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_67_2398 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_67_240 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_67_2406 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_67_2410 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_67_2430 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_67_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_67_2446 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_67_2450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_67_2452 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_67_2469 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_67_2477 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_67_2481 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_67_2484 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_67_2500 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_67_2518 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_67_2522 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_67_2538 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_67_2546 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_67_255 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_67_2562 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_67_2578 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_67_2582 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_67_2586 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_67_2594 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_67_2596 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_67_2609 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_67_2617 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_67_2620 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_67_271 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_67_274 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_67_290 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_67_292 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_67_303 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_67_305 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_67_308 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_67_324 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_67_332 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_67_336 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_67_342 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_67_351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_67_36 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_67_367 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_67_371 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_67_373 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_67_376 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_67_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_67_388 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_67_399 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_67_407 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_67_410 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_67_426 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_67_434 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_67_438 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_67_452 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_67_468 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_67_478 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_67_482 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_67_484 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_67_495 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_67_503 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_67_507 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_67_509 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_67_512 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_67_528 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_67_532 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_67_543 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_67_546 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_67_580 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_67_582 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_67_609 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_67_611 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_67_614 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_67_618 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_67_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_67_642 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_67_648 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_67_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_67_708 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_67_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_67_716 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_67_720 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_67_750 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_67_754 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_67_770 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_67_778 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_67_810 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_67_814 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_67_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_67_822 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_67_849 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_67_852 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_67_856 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_67_86 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_67_872 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_67_880 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_67_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_67_94 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_67_946 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_67_950 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_67_954 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_67_962 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_67_964 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_67_975 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_67_98 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_67_983 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_67_985 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_67_988 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_6_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_6_1011 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_6_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_6_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_6_1081 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_6_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_6_1151 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_6_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_6_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_6_1227 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_6_1291 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_6_1297 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_6_1361 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_6_1367 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_6_1431 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_6_1437 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_6_1501 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_6_1507 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_6_1571 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_6_1577 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_6_1641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_6_1647 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_6_1655 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_6_1659 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_6_1674 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_6_1685 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_6_1689 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_6_1693 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_6_1709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_6_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_6_1713 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_6_1717 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_6_1749 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_6_1757 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_6_1761 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_6_1763 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_6_1766 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_6_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_6_1776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_6_1778 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_6_1821 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_6_1851 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_6_1857 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_6_1859 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_6_1886 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_6_1890 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_6_1894 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_6_1910 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_6_1918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_6_1922 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_6_1924 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_6_1927 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_6_1934 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_6_1950 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_6_1967 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_6_1971 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_6_1987 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_6_1997 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_6_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_6_2061 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_6_2067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_6_2131 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_6_2137 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_6_2201 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_6_2207 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_6_2271 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_6_2277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_6_2341 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_6_2347 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_6_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_6_2411 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_6_2417 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_6_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_6_2481 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_6_2487 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_6_2551 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_6_2557 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_6_2621 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_6_2627 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_6_2643 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_6_2651 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_6_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_6_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_6_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_6_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_6_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_6_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_6_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_6_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_6_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_6_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_6_591 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_6_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_6_661 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_6_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_6_731 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_6_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_6_801 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_6_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_6_871 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_6_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_6_941 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_6_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_7_1046 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_7_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_7_1116 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_7_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_7_1186 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_7_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_7_1256 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_7_1262 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_7_1326 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_7_1332 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_7_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_7_1396 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_7_1402 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_7_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_7_1466 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_7_1472 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_7_1536 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_7_1542 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_7_1606 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_7_1612 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_7_1644 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_7_1660 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_7_1668 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_7_1672 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_7_1676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_7_1682 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_7_1698 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_7_1702 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_7_1736 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_7_1740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_7_1748 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_7_1752 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_7_1792 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_7_1796 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_7_1804 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_7_1808 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_7_1816 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_7_1822 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_7_1832 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_7_1840 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_7_1848 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_7_1900 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_7_1916 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_7_1929 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_7_1946 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_7_1950 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_7_1971 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_7_1975 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_7_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_7_2007 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_7_2023 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_7_2027 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_7_2029 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_7_2032 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_7_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_7_2096 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_7_2102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_7_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_7_2166 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_7_2172 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_7_2236 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_7_2242 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_7_2306 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_7_2312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_7_2376 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_7_2382 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_7_2446 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_7_2452 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_7_2516 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_7_2522 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_7_2586 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_7_2592 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_7_2624 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_7_2640 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_7_2648 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_7_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_7_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_7_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_7_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_7_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_7_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_7_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_7_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_7_556 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_7_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_7_626 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_7_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_7_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_7_696 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_7_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_7_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_7_766 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_7_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_7_836 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_7_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_7_906 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_7_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_7_976 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_7_982 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_8_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_8_1011 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_8_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_8_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_8_1081 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_8_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_8_1151 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_8_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_8_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_8_1227 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_8_1291 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_8_1297 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_8_1361 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_8_1367 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_8_1431 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_8_1437 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_8_1501 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_8_1507 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_8_1571 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_8_1577 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_8_1641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_8_1647 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_8_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_8_1711 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_8_1717 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_8_1749 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_8_1765 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_8_1768 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_8_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_8_1772 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_8_1776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_8_1780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_8_1784 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_8_1787 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_8_1851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_8_1857 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_8_1865 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_8_1869 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_8_1888 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_8_1920 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_8_1924 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_8_1927 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_8_1931 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_8_1947 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_8_1955 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_8_1959 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_8_1962 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_8_1994 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_8_1997 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_8_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_8_2061 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_8_2067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_8_2131 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_8_2137 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_8_2201 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_8_2207 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_8_2271 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_8_2277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_8_2341 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_8_2347 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_8_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_8_2411 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_8_2417 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_8_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_8_2481 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_8_2487 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_8_2551 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_8_2557 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_8_2621 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_8_2627 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_8_2643 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_8_2651 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_8_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_8_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_8_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_8_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_8_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_8_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_8_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_8_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_8_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_8_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_8_591 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_8_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_8_661 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_8_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_8_731 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_8_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_8_801 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_8_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_8_871 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_8_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_8_941 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_8_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_9_1046 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_9_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_9_1116 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_9_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_9_1186 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_9_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_9_1256 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_9_1262 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_9_1326 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_9_1332 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_9_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_9_1396 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_9_1402 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_9_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_9_1466 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_9_1472 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_9_1536 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_9_1542 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_9_1606 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_9_1612 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_9_1676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_9_1682 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_9_1746 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_9_1752 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_9_1816 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_9_1822 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_9_1854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_9_1870 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_9_1878 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_9_1882 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_9_1892 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_9_1956 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_9_1962 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_9_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_9_2026 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_9_2032 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_9_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_9_2096 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_9_2102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_9_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_9_2166 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_9_2172 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_9_2236 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_9_2242 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_9_2306 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_9_2312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_9_2376 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_9_2382 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_9_2446 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_9_2452 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_9_2516 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_9_2522 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_9_2586 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_9_2592 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_9_2624 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_9_2640 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_9_2648 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_9_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_9_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_9_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_9_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_9_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_9_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_9_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_9_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_9_556 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_9_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_9_626 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_9_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_9_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_9_696 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_9_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_9_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_9_766 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_9_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_9_836 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_9_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_9_906 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_9_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_9_976 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_9_982 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_0_Left_68 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_0_Right_0 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_10_Left_78 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_10_Right_10 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_11_Left_79 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_11_Right_11 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_12_Left_80 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_12_Right_12 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_13_Left_81 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_13_Right_13 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_14_Left_82 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_14_Right_14 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_15_Left_83 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_15_Right_15 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_16_Left_84 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_16_Right_16 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_17_Left_85 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_17_Right_17 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_18_Left_86 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_18_Right_18 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_19_Left_87 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_19_Right_19 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_1_Left_69 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_1_Right_1 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_20_Left_88 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_20_Right_20 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_21_Left_89 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_21_Right_21 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_22_Left_90 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_22_Right_22 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_23_Left_91 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_23_Right_23 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_24_Left_92 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_24_Right_24 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_25_Left_93 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_25_Right_25 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_26_Left_94 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_26_Right_26 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_27_Left_95 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_27_Right_27 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_28_Left_96 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_28_Right_28 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_29_Left_97 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_29_Right_29 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_2_Left_70 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_2_Right_2 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_30_Left_98 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_30_Right_30 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_31_Left_99 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_31_Right_31 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_32_Left_100 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_32_Right_32 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_33_Left_101 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_33_Right_33 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_34_Left_102 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_34_Right_34 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_35_Left_103 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_35_Right_35 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_36_Left_104 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_36_Right_36 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_37_Left_105 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_37_Right_37 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_38_Left_106 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_38_Right_38 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_39_Left_107 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_39_Right_39 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_3_Left_71 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_3_Right_3 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_40_Left_108 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_40_Right_40 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_41_Left_109 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_41_Right_41 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_42_Left_110 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_42_Right_42 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_43_Left_111 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_43_Right_43 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_44_Left_112 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_44_Right_44 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_45_Left_113 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_45_Right_45 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_46_Left_114 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_46_Right_46 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_47_Left_115 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_47_Right_47 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_48_Left_116 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_48_Right_48 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_49_Left_117 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_49_Right_49 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_4_Left_72 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_4_Right_4 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_50_Left_118 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_50_Right_50 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_51_Left_119 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_51_Right_51 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_52_Left_120 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_52_Right_52 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_53_Left_121 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_53_Right_53 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_54_Left_122 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_54_Right_54 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_55_Left_123 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_55_Right_55 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_56_Left_124 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_56_Right_56 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_57_Left_125 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_57_Right_57 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_58_Left_126 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_58_Right_58 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_59_Left_127 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_59_Right_59 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_5_Left_73 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_5_Right_5 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_60_Left_128 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_60_Right_60 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_61_Left_129 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_61_Right_61 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_62_Left_130 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_62_Right_62 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_63_Left_131 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_63_Right_63 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_64_Left_132 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_64_Right_64 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_65_Left_133 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_65_Right_65 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_66_Left_134 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_66_Right_66 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_67_Left_135 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_67_Right_67 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_6_Left_74 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_6_Right_6 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_7_Left_75 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_7_Right_7 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_8_Left_76 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_8_Right_8 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_9_Left_77 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_9_Right_9 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_136 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_137 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_138 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_139 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_140 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_141 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_142 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_143 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_144 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_145 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_146 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_147 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_148 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_149 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_150 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_151 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_152 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_153 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_154 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_155 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_156 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_157 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_158 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_159 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_160 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_161 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_162 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_163 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_164 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_165 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_166 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_167 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_168 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_169 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_170 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_171 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_172 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_173 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_174 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_175 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_176 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_177 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_178 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_179 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_180 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_181 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_182 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_183 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_184 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_185 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_186 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_187 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_188 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_189 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_190 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_191 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_192 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_193 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_194 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_195 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_196 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_197 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_198 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_199 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_200 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_201 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_202 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_203 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_204 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_205 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_206 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_207 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_208 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_209 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_210 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_211 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_212 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_10_550 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_10_551 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_10_552 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_10_553 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_10_554 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_10_555 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_10_556 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_10_557 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_10_558 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_10_559 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_10_560 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_10_561 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_10_562 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_10_563 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_10_564 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_10_565 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_10_566 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_10_567 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_10_568 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_10_569 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_10_570 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_10_571 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_10_572 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_10_573 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_10_574 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_10_575 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_10_576 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_10_577 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_10_578 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_10_579 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_10_580 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_10_581 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_10_582 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_10_583 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_10_584 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_10_585 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_10_586 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_10_587 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_11_588 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_11_589 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_11_590 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_11_591 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_11_592 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_11_593 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_11_594 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_11_595 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_11_596 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_11_597 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_11_598 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_11_599 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_11_600 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_11_601 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_11_602 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_11_603 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_11_604 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_11_605 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_11_606 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_11_607 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_11_608 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_11_609 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_11_610 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_11_611 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_11_612 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_11_613 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_11_614 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_11_615 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_11_616 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_11_617 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_11_618 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_11_619 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_11_620 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_11_621 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_11_622 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_11_623 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_11_624 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_12_625 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_12_626 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_12_627 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_12_628 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_12_629 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_12_630 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_12_631 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_12_632 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_12_633 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_12_634 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_12_635 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_12_636 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_12_637 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_12_638 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_12_639 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_12_640 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_12_641 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_12_642 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_12_643 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_12_644 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_12_645 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_12_646 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_12_647 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_12_648 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_12_649 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_12_650 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_12_651 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_12_652 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_12_653 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_12_654 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_12_655 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_12_656 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_12_657 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_12_658 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_12_659 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_12_660 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_12_661 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_12_662 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_13_663 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_13_664 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_13_665 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_13_666 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_13_667 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_13_668 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_13_669 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_13_670 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_13_671 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_13_672 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_13_673 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_13_674 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_13_675 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_13_676 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_13_677 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_13_678 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_13_679 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_13_680 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_13_681 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_13_682 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_13_683 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_13_684 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_13_685 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_13_686 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_13_687 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_13_688 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_13_689 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_13_690 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_13_691 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_13_692 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_13_693 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_13_694 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_13_695 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_13_696 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_13_697 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_13_698 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_13_699 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_14_700 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_14_701 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_14_702 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_14_703 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_14_704 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_14_705 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_14_706 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_14_707 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_14_708 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_14_709 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_14_710 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_14_711 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_14_712 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_14_713 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_14_714 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_14_715 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_14_716 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_14_717 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_14_718 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_14_719 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_14_720 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_14_721 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_14_722 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_14_723 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_14_724 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_14_725 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_14_726 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_14_727 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_14_728 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_14_729 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_14_730 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_14_731 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_14_732 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_14_733 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_14_734 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_14_735 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_14_736 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_14_737 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_15_738 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_15_739 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_15_740 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_15_741 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_15_742 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_15_743 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_15_744 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_15_745 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_15_746 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_15_747 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_15_748 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_15_749 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_15_750 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_15_751 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_15_752 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_15_753 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_15_754 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_15_755 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_15_756 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_15_757 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_15_758 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_15_759 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_15_760 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_15_761 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_15_762 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_15_763 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_15_764 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_15_765 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_15_766 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_15_767 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_15_768 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_15_769 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_15_770 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_15_771 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_15_772 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_15_773 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_15_774 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_16_775 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_16_776 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_16_777 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_16_778 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_16_779 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_16_780 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_16_781 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_16_782 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_16_783 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_16_784 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_16_785 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_16_786 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_16_787 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_16_788 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_16_789 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_16_790 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_16_791 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_16_792 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_16_793 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_16_794 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_16_795 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_16_796 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_16_797 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_16_798 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_16_799 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_16_800 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_16_801 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_16_802 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_16_803 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_16_804 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_16_805 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_16_806 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_16_807 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_16_808 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_16_809 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_16_810 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_16_811 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_16_812 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_17_813 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_17_814 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_17_815 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_17_816 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_17_817 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_17_818 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_17_819 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_17_820 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_17_821 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_17_822 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_17_823 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_17_824 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_17_825 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_17_826 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_17_827 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_17_828 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_17_829 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_17_830 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_17_831 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_17_832 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_17_833 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_17_834 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_17_835 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_17_836 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_17_837 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_17_838 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_17_839 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_17_840 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_17_841 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_17_842 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_17_843 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_17_844 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_17_845 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_17_846 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_17_847 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_17_848 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_17_849 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_18_850 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_18_851 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_18_852 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_18_853 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_18_854 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_18_855 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_18_856 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_18_857 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_18_858 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_18_859 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_18_860 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_18_861 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_18_862 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_18_863 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_18_864 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_18_865 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_18_866 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_18_867 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_18_868 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_18_869 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_18_870 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_18_871 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_18_872 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_18_873 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_18_874 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_18_875 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_18_876 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_18_877 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_18_878 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_18_879 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_18_880 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_18_881 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_18_882 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_18_883 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_18_884 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_18_885 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_18_886 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_18_887 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_19_888 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_19_889 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_19_890 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_19_891 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_19_892 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_19_893 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_19_894 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_19_895 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_19_896 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_19_897 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_19_898 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_19_899 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_19_900 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_19_901 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_19_902 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_19_903 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_19_904 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_19_905 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_19_906 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_19_907 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_19_908 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_19_909 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_19_910 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_19_911 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_19_912 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_19_913 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_19_914 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_19_915 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_19_916 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_19_917 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_19_918 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_19_919 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_19_920 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_19_921 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_19_922 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_19_923 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_19_924 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_1_213 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_1_214 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_1_215 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_1_216 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_1_217 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_1_218 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_1_219 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_1_220 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_1_221 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_1_222 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_1_223 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_1_224 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_1_225 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_1_226 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_1_227 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_1_228 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_1_229 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_1_230 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_1_231 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_1_232 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_1_233 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_1_234 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_1_235 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_1_236 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_1_237 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_1_238 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_1_239 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_1_240 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_1_241 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_1_242 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_1_243 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_1_244 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_1_245 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_1_246 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_1_247 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_1_248 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_1_249 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_20_925 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_20_926 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_20_927 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_20_928 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_20_929 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_20_930 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_20_931 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_20_932 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_20_933 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_20_934 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_20_935 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_20_936 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_20_937 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_20_938 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_20_939 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_20_940 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_20_941 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_20_942 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_20_943 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_20_944 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_20_945 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_20_946 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_20_947 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_20_948 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_20_949 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_20_950 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_20_951 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_20_952 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_20_953 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_20_954 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_20_955 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_20_956 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_20_957 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_20_958 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_20_959 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_20_960 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_20_961 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_20_962 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_21_963 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_21_964 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_21_965 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_21_966 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_21_967 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_21_968 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_21_969 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_21_970 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_21_971 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_21_972 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_21_973 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_21_974 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_21_975 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_21_976 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_21_977 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_21_978 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_21_979 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_21_980 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_21_981 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_21_982 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_21_983 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_21_984 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_21_985 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_21_986 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_21_987 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_21_988 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_21_989 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_21_990 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_21_991 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_21_992 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_21_993 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_21_994 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_21_995 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_21_996 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_21_997 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_21_998 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_21_999 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_22_1000 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_22_1001 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_22_1002 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_22_1003 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_22_1004 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_22_1005 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_22_1006 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_22_1007 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_22_1008 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_22_1009 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_22_1010 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_22_1011 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_22_1012 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_22_1013 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_22_1014 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_22_1015 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_22_1016 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_22_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_22_1018 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_22_1019 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_22_1020 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_22_1021 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_22_1022 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_22_1023 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_22_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_22_1025 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_22_1026 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_22_1027 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_22_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_22_1029 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_22_1030 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_22_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_22_1032 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_22_1033 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_22_1034 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_22_1035 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_22_1036 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_22_1037 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_23_1038 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_23_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_23_1040 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_23_1041 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_23_1042 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_23_1043 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_23_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_23_1045 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_23_1046 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_23_1047 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_23_1048 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_23_1049 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_23_1050 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_23_1051 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_23_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_23_1053 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_23_1054 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_23_1055 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_23_1056 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_23_1057 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_23_1058 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_23_1059 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_23_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_23_1061 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_23_1062 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_23_1063 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_23_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_23_1065 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_23_1066 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_23_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_23_1068 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_23_1069 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_23_1070 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_23_1071 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_23_1072 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_23_1073 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_23_1074 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_24_1075 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_24_1076 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_24_1077 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_24_1078 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_24_1079 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_24_1080 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_24_1081 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_24_1082 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_24_1083 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_24_1084 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_24_1085 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_24_1086 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_24_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_24_1088 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_24_1089 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_24_1090 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_24_1091 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_24_1092 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_24_1093 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_24_1094 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_24_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_24_1096 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_24_1097 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_24_1098 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_24_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_24_1100 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_24_1101 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_24_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_24_1103 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_24_1104 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_24_1105 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_24_1106 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_24_1107 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_24_1108 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_24_1109 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_24_1110 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_24_1111 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_24_1112 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_25_1113 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_25_1114 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_25_1115 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_25_1116 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_25_1117 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_25_1118 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_25_1119 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_25_1120 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_25_1121 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_25_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_25_1123 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_25_1124 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_25_1125 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_25_1126 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_25_1127 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_25_1128 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_25_1129 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_25_1130 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_25_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_25_1132 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_25_1133 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_25_1134 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_25_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_25_1136 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_25_1137 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_25_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_25_1139 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_25_1140 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_25_1141 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_25_1142 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_25_1143 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_25_1144 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_25_1145 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_25_1146 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_25_1147 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_25_1148 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_25_1149 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_26_1150 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_26_1151 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_26_1152 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_26_1153 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_26_1154 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_26_1155 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_26_1156 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_26_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_26_1158 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_26_1159 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_26_1160 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_26_1161 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_26_1162 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_26_1163 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_26_1164 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_26_1165 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_26_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_26_1167 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_26_1168 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_26_1169 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_26_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_26_1171 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_26_1172 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_26_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_26_1174 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_26_1175 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_26_1176 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_26_1177 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_26_1178 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_26_1179 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_26_1180 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_26_1181 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_26_1182 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_26_1183 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_26_1184 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_26_1185 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_26_1186 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_26_1187 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_27_1188 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_27_1189 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_27_1190 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_27_1191 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_27_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_27_1193 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_27_1194 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_27_1195 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_27_1196 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_27_1197 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_27_1198 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_27_1199 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_27_1200 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_27_1201 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_27_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_27_1203 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_27_1204 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_27_1205 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_27_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_27_1207 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_27_1208 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_27_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_27_1210 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_27_1211 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_27_1212 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_27_1213 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_27_1214 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_27_1215 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_27_1216 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_27_1217 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_27_1218 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_27_1219 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_27_1220 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_27_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_27_1222 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_27_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_27_1224 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_28_1225 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_28_1226 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_28_1227 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_28_1228 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_28_1229 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_28_1230 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_28_1231 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_28_1232 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_28_1233 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_28_1234 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_28_1235 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_28_1236 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_28_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_28_1238 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_28_1239 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_28_1240 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_28_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_28_1242 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_28_1243 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_28_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_28_1245 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_28_1246 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_28_1247 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_28_1248 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_28_1249 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_28_1250 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_28_1251 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_28_1252 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_28_1253 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_28_1254 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_28_1255 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_28_1256 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_28_1257 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_28_1258 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_28_1259 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_28_1260 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_28_1261 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_28_1262 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_29_1263 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_29_1264 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_29_1265 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_29_1266 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_29_1267 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_29_1268 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_29_1269 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_29_1270 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_29_1271 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_29_1272 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_29_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_29_1274 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_29_1275 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_29_1276 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_29_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_29_1278 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_29_1279 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_29_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_29_1281 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_29_1282 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_29_1283 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_29_1284 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_29_1285 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_29_1286 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_29_1287 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_29_1288 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_29_1289 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_29_1290 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_29_1291 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_29_1292 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_29_1293 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_29_1294 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_29_1295 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_29_1296 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_29_1297 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_29_1298 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_29_1299 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_2_250 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_2_251 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_2_252 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_2_253 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_2_254 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_2_255 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_2_256 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_2_257 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_2_258 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_2_259 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_2_260 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_2_261 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_2_262 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_2_263 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_2_264 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_2_265 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_2_266 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_2_267 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_2_268 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_2_269 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_2_270 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_2_271 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_2_272 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_2_273 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_2_274 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_2_275 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_2_276 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_2_277 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_2_278 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_2_279 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_2_280 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_2_281 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_2_282 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_2_283 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_2_284 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_2_285 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_2_286 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_2_287 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_30_1300 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_30_1301 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_30_1302 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_30_1303 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_30_1304 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_30_1305 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_30_1306 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_30_1307 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_30_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_30_1309 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_30_1310 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_30_1311 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_30_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_30_1313 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_30_1314 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_30_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_30_1316 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_30_1317 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_30_1318 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_30_1319 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_30_1320 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_30_1321 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_30_1322 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_30_1323 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_30_1324 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_30_1325 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_30_1326 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_30_1327 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_30_1328 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_30_1329 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_30_1330 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_30_1331 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_30_1332 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_30_1333 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_30_1334 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_30_1335 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_30_1336 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_30_1337 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_31_1338 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_31_1339 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_31_1340 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_31_1341 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_31_1342 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_31_1343 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_31_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_31_1345 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_31_1346 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_31_1347 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_31_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_31_1349 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_31_1350 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_31_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_31_1352 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_31_1353 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_31_1354 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_31_1355 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_31_1356 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_31_1357 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_31_1358 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_31_1359 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_31_1360 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_31_1361 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_31_1362 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_31_1363 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_31_1364 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_31_1365 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_31_1366 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_31_1367 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_31_1368 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_31_1369 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_31_1370 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_31_1371 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_31_1372 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_31_1373 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_31_1374 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_32_1375 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_32_1376 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_32_1377 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_32_1378 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_32_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_32_1380 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_32_1381 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_32_1382 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_32_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_32_1384 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_32_1385 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_32_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_32_1387 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_32_1388 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_32_1389 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_32_1390 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_32_1391 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_32_1392 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_32_1393 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_32_1394 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_32_1395 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_32_1396 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_32_1397 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_32_1398 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_32_1399 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_32_1400 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_32_1401 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_32_1402 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_32_1403 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_32_1404 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_32_1405 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_32_1406 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_32_1407 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_32_1408 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_32_1409 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_32_1410 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_32_1411 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_32_1412 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_33_1413 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_33_1414 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_33_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_33_1416 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_33_1417 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_33_1418 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_33_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_33_1420 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_33_1421 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_33_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_33_1423 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_33_1424 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_33_1425 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_33_1426 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_33_1427 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_33_1428 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_33_1429 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_33_1430 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_33_1431 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_33_1432 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_33_1433 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_33_1434 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_33_1435 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_33_1436 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_33_1437 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_33_1438 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_33_1439 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_33_1440 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_33_1441 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_33_1442 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_33_1443 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_33_1444 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_33_1445 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_33_1446 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_33_1447 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_33_1448 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_33_1449 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_34_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_34_1451 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_34_1452 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_34_1453 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_34_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_34_1455 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_34_1456 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_34_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_34_1458 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_34_1459 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_34_1460 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_34_1461 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_34_1462 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_34_1463 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_34_1464 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_34_1465 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_34_1466 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_34_1467 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_34_1468 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_34_1469 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_34_1470 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_34_1471 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_34_1472 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_34_1473 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_34_1474 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_34_1475 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_34_1476 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_34_1477 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_34_1478 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_34_1479 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_34_1480 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_34_1481 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_34_1482 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_34_1483 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_34_1484 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_34_1485 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_34_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_34_1487 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_35_1488 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_35_1489 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_35_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_35_1491 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_35_1492 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_35_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_35_1494 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_35_1495 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_35_1496 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_35_1497 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_35_1498 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_35_1499 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_35_1500 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_35_1501 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_35_1502 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_35_1503 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_35_1504 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_35_1505 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_35_1506 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_35_1507 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_35_1508 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_35_1509 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_35_1510 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_35_1511 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_35_1512 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_35_1513 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_35_1514 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_35_1515 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_35_1516 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_35_1517 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_35_1518 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_35_1519 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_35_1520 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_35_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_35_1522 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_35_1523 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_35_1524 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_36_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_36_1526 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_36_1527 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_36_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_36_1529 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_36_1530 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_36_1531 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_36_1532 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_36_1533 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_36_1534 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_36_1535 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_36_1536 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_36_1537 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_36_1538 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_36_1539 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_36_1540 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_36_1541 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_36_1542 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_36_1543 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_36_1544 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_36_1545 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_36_1546 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_36_1547 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_36_1548 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_36_1549 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_36_1550 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_36_1551 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_36_1552 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_36_1553 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_36_1554 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_36_1555 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_36_1556 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_36_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_36_1558 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_36_1559 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_36_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_36_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_36_1562 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_37_1563 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_37_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_37_1565 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_37_1566 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_37_1567 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_37_1568 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_37_1569 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_37_1570 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_37_1571 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_37_1572 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_37_1573 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_37_1574 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_37_1575 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_37_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_37_1577 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_37_1578 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_37_1579 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_37_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_37_1581 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_37_1582 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_37_1583 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_37_1584 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_37_1585 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_37_1586 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_37_1587 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_37_1588 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_37_1589 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_37_1590 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_37_1591 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_37_1592 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_37_1593 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_37_1594 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_37_1595 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_37_1596 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_37_1597 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_37_1598 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_37_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_38_1600 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_38_1601 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_38_1602 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_38_1603 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_38_1604 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_38_1605 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_38_1606 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_38_1607 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_38_1608 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_38_1609 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_38_1610 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_38_1611 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_38_1612 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_38_1613 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_38_1614 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_38_1615 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_38_1616 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_38_1617 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_38_1618 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_38_1619 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_38_1620 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_38_1621 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_38_1622 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_38_1623 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_38_1624 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_38_1625 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_38_1626 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_38_1627 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_38_1628 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_38_1629 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_38_1630 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_38_1631 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_38_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_38_1633 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_38_1634 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_38_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_38_1636 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_38_1637 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_39_1638 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_39_1639 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_39_1640 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_39_1641 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_39_1642 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_39_1643 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_39_1644 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_39_1645 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_39_1646 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_39_1647 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_39_1648 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_39_1649 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_39_1650 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_39_1651 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_39_1652 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_39_1653 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_39_1654 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_39_1655 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_39_1656 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_39_1657 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_39_1658 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_39_1659 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_39_1660 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_39_1661 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_39_1662 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_39_1663 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_39_1664 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_39_1665 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_39_1666 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_39_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_39_1668 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_39_1669 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_39_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_39_1671 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_39_1672 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_39_1673 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_39_1674 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_3_288 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_3_289 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_3_290 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_3_291 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_3_292 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_3_293 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_3_294 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_3_295 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_3_296 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_3_297 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_3_298 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_3_299 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_3_300 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_3_301 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_3_302 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_3_303 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_3_304 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_3_305 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_3_306 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_3_307 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_3_308 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_3_309 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_3_310 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_3_311 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_3_312 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_3_313 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_3_314 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_3_315 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_3_316 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_3_317 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_3_318 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_3_319 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_3_320 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_3_321 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_3_322 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_3_323 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_3_324 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_40_1675 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_40_1676 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_40_1677 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_40_1678 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_40_1679 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_40_1680 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_40_1681 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_40_1682 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_40_1683 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_40_1684 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_40_1685 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_40_1686 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_40_1687 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_40_1688 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_40_1689 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_40_1690 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_40_1691 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_40_1692 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_40_1693 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_40_1694 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_40_1695 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_40_1696 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_40_1697 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_40_1698 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_40_1699 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_40_1700 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_40_1701 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_40_1702 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_40_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_40_1704 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_40_1705 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_40_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_40_1707 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_40_1708 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_40_1709 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_40_1710 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_40_1711 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_40_1712 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_41_1713 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_41_1714 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_41_1715 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_41_1716 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_41_1717 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_41_1718 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_41_1719 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_41_1720 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_41_1721 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_41_1722 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_41_1723 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_41_1724 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_41_1725 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_41_1726 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_41_1727 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_41_1728 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_41_1729 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_41_1730 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_41_1731 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_41_1732 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_41_1733 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_41_1734 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_41_1735 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_41_1736 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_41_1737 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_41_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_41_1739 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_41_1740 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_41_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_41_1742 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_41_1743 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_41_1744 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_41_1745 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_41_1746 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_41_1747 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_41_1748 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_41_1749 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_42_1750 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_42_1751 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_42_1752 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_42_1753 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_42_1754 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_42_1755 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_42_1756 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_42_1757 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_42_1758 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_42_1759 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_42_1760 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_42_1761 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_42_1762 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_42_1763 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_42_1764 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_42_1765 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_42_1766 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_42_1767 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_42_1768 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_42_1769 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_42_1770 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_42_1771 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_42_1772 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_42_1773 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_42_1774 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_42_1775 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_42_1776 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_42_1777 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_42_1778 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_42_1779 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_42_1780 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_42_1781 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_42_1782 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_42_1783 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_42_1784 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_42_1785 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_42_1786 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_42_1787 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_43_1788 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_43_1789 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_43_1790 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_43_1791 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_43_1792 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_43_1793 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_43_1794 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_43_1795 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_43_1796 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_43_1797 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_43_1798 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_43_1799 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_43_1800 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_43_1801 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_43_1802 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_43_1803 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_43_1804 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_43_1805 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_43_1806 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_43_1807 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_43_1808 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_43_1809 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_43_1810 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_43_1811 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_43_1812 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_43_1813 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_43_1814 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_43_1815 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_43_1816 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_43_1817 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_43_1818 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_43_1819 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_43_1820 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_43_1821 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_43_1822 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_43_1823 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_43_1824 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_44_1825 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_44_1826 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_44_1827 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_44_1828 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_44_1829 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_44_1830 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_44_1831 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_44_1832 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_44_1833 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_44_1834 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_44_1835 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_44_1836 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_44_1837 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_44_1838 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_44_1839 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_44_1840 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_44_1841 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_44_1842 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_44_1843 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_44_1844 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_44_1845 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_44_1846 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_44_1847 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_44_1848 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_44_1849 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_44_1850 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_44_1851 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_44_1852 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_44_1853 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_44_1854 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_44_1855 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_44_1856 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_44_1857 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_44_1858 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_44_1859 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_44_1860 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_44_1861 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_44_1862 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_45_1863 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_45_1864 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_45_1865 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_45_1866 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_45_1867 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_45_1868 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_45_1869 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_45_1870 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_45_1871 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_45_1872 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_45_1873 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_45_1874 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_45_1875 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_45_1876 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_45_1877 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_45_1878 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_45_1879 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_45_1880 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_45_1881 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_45_1882 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_45_1883 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_45_1884 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_45_1885 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_45_1886 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_45_1887 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_45_1888 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_45_1889 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_45_1890 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_45_1891 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_45_1892 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_45_1893 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_45_1894 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_45_1895 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_45_1896 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_45_1897 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_45_1898 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_45_1899 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_46_1900 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_46_1901 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_46_1902 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_46_1903 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_46_1904 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_46_1905 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_46_1906 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_46_1907 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_46_1908 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_46_1909 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_46_1910 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_46_1911 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_46_1912 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_46_1913 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_46_1914 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_46_1915 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_46_1916 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_46_1917 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_46_1918 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_46_1919 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_46_1920 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_46_1921 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_46_1922 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_46_1923 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_46_1924 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_46_1925 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_46_1926 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_46_1927 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_46_1928 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_46_1929 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_46_1930 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_46_1931 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_46_1932 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_46_1933 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_46_1934 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_46_1935 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_46_1936 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_46_1937 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_47_1938 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_47_1939 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_47_1940 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_47_1941 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_47_1942 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_47_1943 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_47_1944 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_47_1945 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_47_1946 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_47_1947 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_47_1948 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_47_1949 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_47_1950 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_47_1951 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_47_1952 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_47_1953 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_47_1954 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_47_1955 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_47_1956 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_47_1957 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_47_1958 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_47_1959 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_47_1960 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_47_1961 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_47_1962 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_47_1963 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_47_1964 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_47_1965 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_47_1966 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_47_1967 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_47_1968 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_47_1969 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_47_1970 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_47_1971 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_47_1972 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_47_1973 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_47_1974 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_48_1975 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_48_1976 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_48_1977 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_48_1978 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_48_1979 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_48_1980 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_48_1981 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_48_1982 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_48_1983 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_48_1984 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_48_1985 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_48_1986 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_48_1987 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_48_1988 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_48_1989 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_48_1990 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_48_1991 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_48_1992 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_48_1993 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_48_1994 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_48_1995 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_48_1996 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_48_1997 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_48_1998 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_48_1999 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_48_2000 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_48_2001 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_48_2002 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_48_2003 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_48_2004 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_48_2005 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_48_2006 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_48_2007 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_48_2008 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_48_2009 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_48_2010 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_48_2011 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_48_2012 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_49_2013 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_49_2014 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_49_2015 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_49_2016 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_49_2017 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_49_2018 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_49_2019 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_49_2020 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_49_2021 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_49_2022 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_49_2023 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_49_2024 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_49_2025 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_49_2026 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_49_2027 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_49_2028 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_49_2029 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_49_2030 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_49_2031 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_49_2032 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_49_2033 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_49_2034 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_49_2035 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_49_2036 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_49_2037 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_49_2038 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_49_2039 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_49_2040 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_49_2041 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_49_2042 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_49_2043 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_49_2044 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_49_2045 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_49_2046 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_49_2047 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_49_2048 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_49_2049 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_4_325 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_4_326 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_4_327 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_4_328 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_4_329 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_4_330 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_4_331 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_4_332 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_4_333 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_4_334 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_4_335 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_4_336 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_4_337 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_4_338 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_4_339 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_4_340 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_4_341 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_4_342 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_4_343 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_4_344 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_4_345 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_4_346 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_4_347 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_4_348 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_4_349 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_4_350 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_4_351 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_4_352 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_4_353 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_4_354 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_4_355 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_4_356 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_4_357 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_4_358 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_4_359 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_4_360 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_4_361 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_4_362 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_50_2050 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_50_2051 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_50_2052 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_50_2053 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_50_2054 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_50_2055 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_50_2056 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_50_2057 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_50_2058 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_50_2059 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_50_2060 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_50_2061 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_50_2062 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_50_2063 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_50_2064 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_50_2065 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_50_2066 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_50_2067 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_50_2068 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_50_2069 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_50_2070 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_50_2071 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_50_2072 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_50_2073 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_50_2074 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_50_2075 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_50_2076 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_50_2077 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_50_2078 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_50_2079 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_50_2080 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_50_2081 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_50_2082 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_50_2083 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_50_2084 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_50_2085 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_50_2086 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_50_2087 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_51_2088 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_51_2089 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_51_2090 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_51_2091 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_51_2092 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_51_2093 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_51_2094 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_51_2095 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_51_2096 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_51_2097 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_51_2098 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_51_2099 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_51_2100 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_51_2101 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_51_2102 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_51_2103 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_51_2104 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_51_2105 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_51_2106 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_51_2107 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_51_2108 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_51_2109 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_51_2110 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_51_2111 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_51_2112 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_51_2113 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_51_2114 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_51_2115 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_51_2116 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_51_2117 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_51_2118 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_51_2119 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_51_2120 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_51_2121 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_51_2122 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_51_2123 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_51_2124 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_52_2125 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_52_2126 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_52_2127 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_52_2128 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_52_2129 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_52_2130 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_52_2131 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_52_2132 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_52_2133 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_52_2134 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_52_2135 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_52_2136 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_52_2137 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_52_2138 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_52_2139 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_52_2140 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_52_2141 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_52_2142 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_52_2143 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_52_2144 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_52_2145 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_52_2146 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_52_2147 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_52_2148 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_52_2149 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_52_2150 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_52_2151 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_52_2152 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_52_2153 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_52_2154 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_52_2155 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_52_2156 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_52_2157 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_52_2158 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_52_2159 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_52_2160 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_52_2161 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_52_2162 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_53_2163 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_53_2164 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_53_2165 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_53_2166 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_53_2167 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_53_2168 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_53_2169 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_53_2170 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_53_2171 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_53_2172 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_53_2173 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_53_2174 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_53_2175 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_53_2176 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_53_2177 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_53_2178 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_53_2179 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_53_2180 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_53_2181 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_53_2182 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_53_2183 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_53_2184 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_53_2185 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_53_2186 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_53_2187 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_53_2188 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_53_2189 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_53_2190 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_53_2191 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_53_2192 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_53_2193 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_53_2194 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_53_2195 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_53_2196 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_53_2197 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_53_2198 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_53_2199 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_54_2200 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_54_2201 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_54_2202 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_54_2203 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_54_2204 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_54_2205 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_54_2206 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_54_2207 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_54_2208 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_54_2209 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_54_2210 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_54_2211 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_54_2212 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_54_2213 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_54_2214 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_54_2215 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_54_2216 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_54_2217 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_54_2218 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_54_2219 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_54_2220 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_54_2221 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_54_2222 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_54_2223 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_54_2224 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_54_2225 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_54_2226 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_54_2227 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_54_2228 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_54_2229 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_54_2230 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_54_2231 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_54_2232 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_54_2233 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_54_2234 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_54_2235 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_54_2236 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_54_2237 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_55_2238 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_55_2239 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_55_2240 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_55_2241 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_55_2242 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_55_2243 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_55_2244 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_55_2245 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_55_2246 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_55_2247 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_55_2248 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_55_2249 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_55_2250 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_55_2251 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_55_2252 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_55_2253 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_55_2254 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_55_2255 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_55_2256 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_55_2257 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_55_2258 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_55_2259 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_55_2260 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_55_2261 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_55_2262 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_55_2263 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_55_2264 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_55_2265 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_55_2266 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_55_2267 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_55_2268 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_55_2269 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_55_2270 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_55_2271 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_55_2272 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_55_2273 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_55_2274 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_56_2275 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_56_2276 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_56_2277 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_56_2278 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_56_2279 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_56_2280 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_56_2281 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_56_2282 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_56_2283 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_56_2284 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_56_2285 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_56_2286 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_56_2287 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_56_2288 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_56_2289 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_56_2290 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_56_2291 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_56_2292 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_56_2293 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_56_2294 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_56_2295 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_56_2296 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_56_2297 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_56_2298 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_56_2299 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_56_2300 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_56_2301 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_56_2302 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_56_2303 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_56_2304 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_56_2305 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_56_2306 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_56_2307 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_56_2308 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_56_2309 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_56_2310 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_56_2311 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_56_2312 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_57_2313 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_57_2314 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_57_2315 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_57_2316 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_57_2317 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_57_2318 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_57_2319 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_57_2320 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_57_2321 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_57_2322 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_57_2323 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_57_2324 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_57_2325 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_57_2326 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_57_2327 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_57_2328 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_57_2329 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_57_2330 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_57_2331 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_57_2332 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_57_2333 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_57_2334 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_57_2335 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_57_2336 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_57_2337 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_57_2338 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_57_2339 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_57_2340 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_57_2341 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_57_2342 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_57_2343 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_57_2344 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_57_2345 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_57_2346 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_57_2347 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_57_2348 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_57_2349 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_58_2350 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_58_2351 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_58_2352 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_58_2353 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_58_2354 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_58_2355 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_58_2356 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_58_2357 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_58_2358 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_58_2359 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_58_2360 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_58_2361 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_58_2362 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_58_2363 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_58_2364 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_58_2365 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_58_2366 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_58_2367 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_58_2368 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_58_2369 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_58_2370 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_58_2371 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_58_2372 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_58_2373 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_58_2374 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_58_2375 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_58_2376 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_58_2377 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_58_2378 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_58_2379 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_58_2380 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_58_2381 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_58_2382 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_58_2383 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_58_2384 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_58_2385 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_58_2386 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_58_2387 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_59_2388 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_59_2389 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_59_2390 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_59_2391 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_59_2392 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_59_2393 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_59_2394 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_59_2395 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_59_2396 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_59_2397 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_59_2398 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_59_2399 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_59_2400 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_59_2401 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_59_2402 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_59_2403 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_59_2404 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_59_2405 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_59_2406 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_59_2407 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_59_2408 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_59_2409 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_59_2410 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_59_2411 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_59_2412 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_59_2413 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_59_2414 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_59_2415 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_59_2416 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_59_2417 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_59_2418 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_59_2419 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_59_2420 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_59_2421 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_59_2422 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_59_2423 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_59_2424 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_5_363 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_5_364 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_5_365 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_5_366 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_5_367 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_5_368 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_5_369 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_5_370 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_5_371 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_5_372 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_5_373 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_5_374 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_5_375 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_5_376 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_5_377 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_5_378 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_5_379 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_5_380 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_5_381 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_5_382 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_5_383 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_5_384 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_5_385 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_5_386 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_5_387 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_5_388 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_5_389 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_5_390 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_5_391 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_5_392 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_5_393 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_5_394 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_5_395 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_5_396 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_5_397 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_5_398 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_5_399 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_60_2425 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_60_2426 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_60_2427 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_60_2428 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_60_2429 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_60_2430 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_60_2431 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_60_2432 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_60_2433 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_60_2434 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_60_2435 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_60_2436 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_60_2437 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_60_2438 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_60_2439 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_60_2440 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_60_2441 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_60_2442 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_60_2443 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_60_2444 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_60_2445 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_60_2446 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_60_2447 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_60_2448 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_60_2449 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_60_2450 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_60_2451 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_60_2452 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_60_2453 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_60_2454 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_60_2455 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_60_2456 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_60_2457 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_60_2458 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_60_2459 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_60_2460 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_60_2461 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_60_2462 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_61_2463 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_61_2464 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_61_2465 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_61_2466 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_61_2467 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_61_2468 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_61_2469 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_61_2470 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_61_2471 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_61_2472 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_61_2473 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_61_2474 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_61_2475 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_61_2476 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_61_2477 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_61_2478 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_61_2479 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_61_2480 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_61_2481 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_61_2482 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_61_2483 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_61_2484 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_61_2485 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_61_2486 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_61_2487 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_61_2488 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_61_2489 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_61_2490 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_61_2491 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_61_2492 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_61_2493 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_61_2494 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_61_2495 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_61_2496 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_61_2497 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_61_2498 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_61_2499 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_62_2500 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_62_2501 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_62_2502 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_62_2503 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_62_2504 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_62_2505 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_62_2506 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_62_2507 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_62_2508 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_62_2509 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_62_2510 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_62_2511 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_62_2512 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_62_2513 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_62_2514 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_62_2515 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_62_2516 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_62_2517 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_62_2518 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_62_2519 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_62_2520 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_62_2521 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_62_2522 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_62_2523 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_62_2524 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_62_2525 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_62_2526 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_62_2527 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_62_2528 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_62_2529 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_62_2530 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_62_2531 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_62_2532 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_62_2533 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_62_2534 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_62_2535 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_62_2536 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_62_2537 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_63_2538 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_63_2539 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_63_2540 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_63_2541 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_63_2542 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_63_2543 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_63_2544 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_63_2545 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_63_2546 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_63_2547 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_63_2548 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_63_2549 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_63_2550 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_63_2551 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_63_2552 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_63_2553 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_63_2554 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_63_2555 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_63_2556 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_63_2557 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_63_2558 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_63_2559 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_63_2560 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_63_2561 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_63_2562 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_63_2563 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_63_2564 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_63_2565 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_63_2566 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_63_2567 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_63_2568 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_63_2569 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_63_2570 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_63_2571 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_63_2572 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_63_2573 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_63_2574 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_64_2575 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_64_2576 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_64_2577 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_64_2578 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_64_2579 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_64_2580 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_64_2581 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_64_2582 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_64_2583 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_64_2584 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_64_2585 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_64_2586 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_64_2587 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_64_2588 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_64_2589 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_64_2590 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_64_2591 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_64_2592 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_64_2593 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_64_2594 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_64_2595 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_64_2596 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_64_2597 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_64_2598 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_64_2599 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_64_2600 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_64_2601 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_64_2602 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_64_2603 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_64_2604 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_64_2605 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_64_2606 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_64_2607 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_64_2608 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_64_2609 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_64_2610 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_64_2611 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_64_2612 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_65_2613 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_65_2614 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_65_2615 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_65_2616 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_65_2617 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_65_2618 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_65_2619 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_65_2620 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_65_2621 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_65_2622 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_65_2623 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_65_2624 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_65_2625 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_65_2626 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_65_2627 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_65_2628 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_65_2629 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_65_2630 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_65_2631 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_65_2632 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_65_2633 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_65_2634 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_65_2635 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_65_2636 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_65_2637 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_65_2638 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_65_2639 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_65_2640 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_65_2641 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_65_2642 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_65_2643 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_65_2644 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_65_2645 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_65_2646 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_65_2647 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_65_2648 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_65_2649 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_66_2650 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_66_2651 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_66_2652 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_66_2653 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_66_2654 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_66_2655 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_66_2656 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_66_2657 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_66_2658 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_66_2659 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_66_2660 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_66_2661 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_66_2662 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_66_2663 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_66_2664 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_66_2665 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_66_2666 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_66_2667 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_66_2668 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_66_2669 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_66_2670 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_66_2671 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_66_2672 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_66_2673 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_66_2674 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_66_2675 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_66_2676 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_66_2677 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_66_2678 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_66_2679 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_66_2680 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_66_2681 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_66_2682 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_66_2683 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_66_2684 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_66_2685 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_66_2686 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_66_2687 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_67_2688 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_67_2689 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_67_2690 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_67_2691 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_67_2692 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_67_2693 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_67_2694 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_67_2695 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_67_2696 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_67_2697 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_67_2698 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_67_2699 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_67_2700 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_67_2701 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_67_2702 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_67_2703 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_67_2704 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_67_2705 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_67_2706 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_67_2707 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_67_2708 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_67_2709 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_67_2710 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_67_2711 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_67_2712 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_67_2713 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_67_2714 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_67_2715 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_67_2716 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_67_2717 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_67_2718 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_67_2719 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_67_2720 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_67_2721 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_67_2722 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_67_2723 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_67_2724 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_67_2725 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_67_2726 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_67_2727 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_67_2728 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_67_2729 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_67_2730 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_67_2731 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_67_2732 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_67_2733 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_67_2734 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_67_2735 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_67_2736 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_67_2737 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_67_2738 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_67_2739 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_67_2740 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_67_2741 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_67_2742 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_67_2743 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_67_2744 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_67_2745 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_67_2746 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_67_2747 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_67_2748 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_67_2749 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_67_2750 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_67_2751 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_67_2752 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_67_2753 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_67_2754 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_67_2755 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_67_2756 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_67_2757 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_67_2758 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_67_2759 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_67_2760 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_67_2761 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_67_2762 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_67_2763 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_67_2764 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_6_400 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_6_401 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_6_402 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_6_403 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_6_404 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_6_405 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_6_406 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_6_407 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_6_408 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_6_409 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_6_410 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_6_411 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_6_412 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_6_413 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_6_414 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_6_415 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_6_416 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_6_417 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_6_418 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_6_419 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_6_420 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_6_421 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_6_422 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_6_423 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_6_424 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_6_425 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_6_426 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_6_427 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_6_428 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_6_429 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_6_430 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_6_431 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_6_432 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_6_433 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_6_434 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_6_435 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_6_436 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_6_437 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_7_438 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_7_439 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_7_440 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_7_441 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_7_442 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_7_443 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_7_444 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_7_445 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_7_446 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_7_447 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_7_448 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_7_449 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_7_450 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_7_451 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_7_452 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_7_453 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_7_454 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_7_455 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_7_456 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_7_457 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_7_458 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_7_459 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_7_460 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_7_461 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_7_462 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_7_463 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_7_464 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_7_465 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_7_466 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_7_467 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_7_468 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_7_469 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_7_470 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_7_471 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_7_472 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_7_473 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_7_474 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_8_475 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_8_476 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_8_477 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_8_478 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_8_479 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_8_480 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_8_481 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_8_482 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_8_483 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_8_484 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_8_485 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_8_486 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_8_487 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_8_488 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_8_489 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_8_490 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_8_491 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_8_492 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_8_493 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_8_494 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_8_495 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_8_496 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_8_497 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_8_498 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_8_499 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_8_500 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_8_501 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_8_502 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_8_503 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_8_504 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_8_505 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_8_506 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_8_507 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_8_508 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_8_509 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_8_510 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_8_511 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_8_512 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_9_513 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_9_514 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_9_515 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_9_516 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_9_517 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_9_518 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_9_519 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_9_520 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_9_521 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_9_522 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_9_523 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_9_524 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_9_525 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_9_526 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_9_527 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_9_528 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_9_529 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_9_530 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_9_531 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_9_532 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_9_533 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_9_534 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_9_535 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_9_536 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_9_537 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_9_538 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_9_539 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_9_540 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_9_541 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_9_542 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_9_543 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_9_544 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_9_545 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_9_546 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_9_547 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_9_548 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_9_549 ();
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _106_ (.I(_004_),
    .Z(_073_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _107_ (.I(_025_),
    .Z(_074_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _108_ (.A1(_073_),
    .A2(_074_),
    .A3(_057_),
    .A4(net52),
    .ZN(_075_));
 gf180mcu_fd_sc_mcu7t5v0__and4_1 _109_ (.A1(_068_),
    .A2(_070_),
    .A3(_072_),
    .A4(_075_),
    .Z(_076_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_4 _110_ (.A1(_060_),
    .A2(_061_),
    .B1(_065_),
    .B2(_076_),
    .ZN(net121));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _111_ (.I(net5),
    .ZN(_077_));
 gf180mcu_fd_sc_mcu7t5v0__aoi222_4 _112_ (.A1(net21),
    .A2(_062_),
    .B1(_063_),
    .B2(net45),
    .C1(net61),
    .C2(_064_),
    .ZN(_078_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_2 _113_ (.A1(_066_),
    .A2(_067_),
    .A3(_051_),
    .A4(net13),
    .ZN(_079_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _114_ (.A1(_053_),
    .A2(net29),
    .A3(_069_),
    .ZN(_080_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _115_ (.A1(_055_),
    .A2(net37),
    .B(_071_),
    .ZN(_081_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _116_ (.A1(_073_),
    .A2(_074_),
    .A3(_057_),
    .A4(net53),
    .ZN(_082_));
 gf180mcu_fd_sc_mcu7t5v0__and4_1 _117_ (.A1(_079_),
    .A2(_080_),
    .A3(_081_),
    .A4(_082_),
    .Z(_083_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_4 _118_ (.A1(_077_),
    .A2(_061_),
    .B1(_078_),
    .B2(_083_),
    .ZN(net122));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _119_ (.I(net6),
    .ZN(_084_));
 gf180mcu_fd_sc_mcu7t5v0__aoi222_4 _120_ (.A1(net22),
    .A2(_062_),
    .B1(_063_),
    .B2(net46),
    .C1(net62),
    .C2(_064_),
    .ZN(_085_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_2 _121_ (.A1(_066_),
    .A2(_067_),
    .A3(_051_),
    .A4(net14),
    .ZN(_086_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _122_ (.A1(_053_),
    .A2(net30),
    .A3(_069_),
    .ZN(_087_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _123_ (.A1(_055_),
    .A2(net38),
    .B(_071_),
    .ZN(_088_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _124_ (.A1(_073_),
    .A2(_074_),
    .A3(_057_),
    .A4(net54),
    .ZN(_089_));
 gf180mcu_fd_sc_mcu7t5v0__and4_1 _125_ (.A1(_086_),
    .A2(_087_),
    .A3(_088_),
    .A4(_089_),
    .Z(_090_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_4 _126_ (.A1(_084_),
    .A2(_061_),
    .B1(_085_),
    .B2(_090_),
    .ZN(net123));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _127_ (.I(net7),
    .ZN(_091_));
 gf180mcu_fd_sc_mcu7t5v0__aoi222_4 _128_ (.A1(net23),
    .A2(_062_),
    .B1(_063_),
    .B2(net47),
    .C1(net63),
    .C2(_064_),
    .ZN(_092_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _129_ (.A1(_066_),
    .A2(_067_),
    .A3(_015_),
    .A4(net15),
    .ZN(_093_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _130_ (.A1(_038_),
    .A2(net31),
    .A3(_069_),
    .ZN(_094_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _131_ (.A1(_035_),
    .A2(net39),
    .B(_071_),
    .ZN(_095_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _132_ (.A1(_073_),
    .A2(_074_),
    .A3(_008_),
    .A4(net55),
    .ZN(_096_));
 gf180mcu_fd_sc_mcu7t5v0__and4_1 _133_ (.A1(_093_),
    .A2(_094_),
    .A3(_095_),
    .A4(_096_),
    .Z(_097_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_4 _134_ (.A1(_091_),
    .A2(_061_),
    .B1(_092_),
    .B2(_097_),
    .ZN(net124));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _135_ (.I(net8),
    .ZN(_098_));
 gf180mcu_fd_sc_mcu7t5v0__aoi222_4 _136_ (.A1(net24),
    .A2(_018_),
    .B1(_026_),
    .B2(net48),
    .C1(net64),
    .C2(_030_),
    .ZN(_099_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _137_ (.A1(_011_),
    .A2(_006_),
    .A3(_015_),
    .A4(net16),
    .ZN(_100_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _138_ (.A1(_038_),
    .A2(net32),
    .A3(_020_),
    .ZN(_101_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _139_ (.A1(_035_),
    .A2(net40),
    .B(_023_),
    .ZN(_102_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _140_ (.A1(_004_),
    .A2(_025_),
    .A3(_008_),
    .A4(net56),
    .ZN(_103_));
 gf180mcu_fd_sc_mcu7t5v0__and4_1 _141_ (.A1(_100_),
    .A2(_101_),
    .A3(_102_),
    .A4(_103_),
    .Z(_104_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_4 _142_ (.A1(_098_),
    .A2(_009_),
    .B1(_099_),
    .B2(_104_),
    .ZN(net125));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _143_ (.A1(\aaaa[14] ),
    .A2(\aaaa[12] ),
    .A3(\aaaa[13] ),
    .ZN(_105_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _144_ (.A1(net74),
    .A2(_105_),
    .ZN(_000_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_4 _145_ (.A1(net65),
    .A2(\aaaa[15] ),
    .A3(_000_),
    .ZN(_001_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _146_ (.I(_001_),
    .Z(_002_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _147_ (.I(\aaaa[1] ),
    .Z(_003_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _148_ (.I(_003_),
    .Z(_004_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _149_ (.I(\aaaa[0] ),
    .Z(_005_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _150_ (.I(_005_),
    .Z(_006_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _151_ (.I(\aaaa[2] ),
    .Z(_007_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _152_ (.I(_007_),
    .Z(_008_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_4 _153_ (.A1(_004_),
    .A2(_006_),
    .A3(_008_),
    .ZN(_009_));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _154_ (.I(_009_),
    .Z(_010_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_4 _155_ (.A1(_002_),
    .A2(_010_),
    .ZN(net110));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _156_ (.I(_003_),
    .ZN(_011_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _157_ (.I(_011_),
    .Z(_012_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _158_ (.I(_006_),
    .Z(_013_));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _159_ (.I(\aaaa[2] ),
    .ZN(_014_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _160_ (.I(_014_),
    .Z(_015_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _161_ (.I(_015_),
    .Z(_016_));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _162_ (.I(_001_),
    .Z(_017_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_4 _163_ (.A1(_012_),
    .A2(_013_),
    .A3(_016_),
    .A4(_017_),
    .ZN(net111));
 gf180mcu_fd_sc_mcu7t5v0__nor3_4 _164_ (.A1(_011_),
    .A2(_005_),
    .A3(_007_),
    .ZN(_018_));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _165_ (.I(_018_),
    .Z(_019_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_4 _166_ (.A1(_002_),
    .A2(_019_),
    .ZN(net112));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _167_ (.A1(\aaaa[1] ),
    .A2(\aaaa[0] ),
    .Z(_020_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _168_ (.I(_020_),
    .Z(_021_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_4 _169_ (.A1(_016_),
    .A2(_017_),
    .A3(_021_),
    .ZN(net113));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _170_ (.I(_008_),
    .Z(_022_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _171_ (.A1(_003_),
    .A2(_005_),
    .ZN(_023_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _172_ (.I(_023_),
    .Z(_024_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_4 _173_ (.A1(_022_),
    .A2(_017_),
    .A3(_024_),
    .ZN(net114));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _174_ (.I(_005_),
    .ZN(_025_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_4 _175_ (.A1(_003_),
    .A2(_025_),
    .A3(_014_),
    .ZN(_026_));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _176_ (.I(_026_),
    .Z(_027_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _177_ (.A1(_002_),
    .A2(_027_),
    .ZN(net115));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _178_ (.I(_004_),
    .Z(_028_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _179_ (.I(_025_),
    .Z(_029_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_4 _180_ (.A1(_028_),
    .A2(_029_),
    .A3(_022_),
    .A4(_017_),
    .ZN(net116));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _181_ (.A1(_007_),
    .A2(_020_),
    .Z(_030_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _182_ (.I(_030_),
    .Z(_031_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _183_ (.A1(_002_),
    .A2(_031_),
    .ZN(net117));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _184_ (.I(net1),
    .ZN(_032_));
 gf180mcu_fd_sc_mcu7t5v0__aoi222_4 _185_ (.A1(net17),
    .A2(_019_),
    .B1(_027_),
    .B2(net41),
    .C1(net57),
    .C2(_031_),
    .ZN(_033_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _186_ (.I(_014_),
    .Z(_034_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _187_ (.I(_034_),
    .Z(_035_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _188_ (.A1(_012_),
    .A2(_013_),
    .A3(_035_),
    .A4(net9),
    .ZN(_036_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _189_ (.A1(_016_),
    .A2(net25),
    .A3(_021_),
    .ZN(_037_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _190_ (.I(_034_),
    .Z(_038_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _191_ (.A1(_038_),
    .A2(net33),
    .B(_024_),
    .ZN(_039_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _192_ (.A1(_028_),
    .A2(_029_),
    .A3(_022_),
    .A4(net49),
    .ZN(_040_));
 gf180mcu_fd_sc_mcu7t5v0__and4_1 _193_ (.A1(_036_),
    .A2(_037_),
    .A3(_039_),
    .A4(_040_),
    .Z(_041_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_4 _194_ (.A1(_032_),
    .A2(_010_),
    .B1(_033_),
    .B2(_041_),
    .ZN(net118));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _195_ (.I(net2),
    .ZN(_042_));
 gf180mcu_fd_sc_mcu7t5v0__aoi222_4 _196_ (.A1(net18),
    .A2(_019_),
    .B1(_027_),
    .B2(net42),
    .C1(net58),
    .C2(_031_),
    .ZN(_043_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _197_ (.A1(_012_),
    .A2(_013_),
    .A3(_035_),
    .A4(net10),
    .ZN(_044_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _198_ (.A1(_016_),
    .A2(net26),
    .A3(_021_),
    .ZN(_045_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _199_ (.A1(_038_),
    .A2(net34),
    .B(_024_),
    .ZN(_046_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _200_ (.A1(_028_),
    .A2(_029_),
    .A3(_022_),
    .A4(net50),
    .ZN(_047_));
 gf180mcu_fd_sc_mcu7t5v0__and4_1 _201_ (.A1(_044_),
    .A2(_045_),
    .A3(_046_),
    .A4(_047_),
    .Z(_048_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_4 _202_ (.A1(_042_),
    .A2(_010_),
    .B1(_043_),
    .B2(_048_),
    .ZN(net119));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _203_ (.I(net3),
    .ZN(_049_));
 gf180mcu_fd_sc_mcu7t5v0__aoi222_4 _204_ (.A1(net19),
    .A2(_019_),
    .B1(_027_),
    .B2(net43),
    .C1(net59),
    .C2(_031_),
    .ZN(_050_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _205_ (.I(_034_),
    .Z(_051_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _206_ (.A1(_012_),
    .A2(_013_),
    .A3(_051_),
    .A4(net11),
    .ZN(_052_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _207_ (.I(_015_),
    .Z(_053_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _208_ (.A1(_053_),
    .A2(net27),
    .A3(_021_),
    .ZN(_054_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _209_ (.I(_034_),
    .Z(_055_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _210_ (.A1(_055_),
    .A2(net35),
    .B(_024_),
    .ZN(_056_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _211_ (.I(_007_),
    .Z(_057_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _212_ (.A1(_028_),
    .A2(_029_),
    .A3(_057_),
    .A4(net51),
    .ZN(_058_));
 gf180mcu_fd_sc_mcu7t5v0__and4_2 _213_ (.A1(_052_),
    .A2(_054_),
    .A3(_056_),
    .A4(_058_),
    .Z(_059_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_4 _214_ (.A1(_049_),
    .A2(_010_),
    .B1(_050_),
    .B2(_059_),
    .ZN(net120));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _215_ (.I(net4),
    .ZN(_060_));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _216_ (.I(_009_),
    .Z(_061_));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _217_ (.I(_018_),
    .Z(_062_));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _218_ (.I(_026_),
    .Z(_063_));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _219_ (.I(_030_),
    .Z(_064_));
 gf180mcu_fd_sc_mcu7t5v0__aoi222_4 _220_ (.A1(net20),
    .A2(_062_),
    .B1(_063_),
    .B2(net44),
    .C1(net60),
    .C2(_064_),
    .ZN(_065_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _221_ (.I(_011_),
    .Z(_066_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _222_ (.I(_006_),
    .Z(_067_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_2 _223_ (.A1(_066_),
    .A2(_067_),
    .A3(_051_),
    .A4(net12),
    .ZN(_068_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _224_ (.I(_020_),
    .Z(_069_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _225_ (.A1(_053_),
    .A2(net28),
    .A3(_069_),
    .ZN(_070_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _226_ (.I(_023_),
    .Z(_071_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _227_ (.A1(_055_),
    .A2(net36),
    .B(_071_),
    .ZN(_072_));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _228_ (.D(net75),
    .CLK(clknet_1_1__leaf_wb_clk_i),
    .Q(\aaaa[0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _229_ (.D(net82),
    .CLK(clknet_1_1__leaf_wb_clk_i),
    .Q(\aaaa[1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _230_ (.D(net83),
    .CLK(clknet_1_1__leaf_wb_clk_i),
    .Q(\aaaa[2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _231_ (.D(net84),
    .CLK(clknet_1_0__leaf_wb_clk_i),
    .Q(\aaaa[3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _232_ (.D(net85),
    .CLK(clknet_1_0__leaf_wb_clk_i),
    .Q(\aaaa[4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _233_ (.D(net86),
    .CLK(clknet_1_0__leaf_wb_clk_i),
    .Q(\aaaa[5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _234_ (.D(net87),
    .CLK(clknet_1_0__leaf_wb_clk_i),
    .Q(\aaaa[6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _235_ (.D(net88),
    .CLK(clknet_1_0__leaf_wb_clk_i),
    .Q(\aaaa[7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _236_ (.D(net89),
    .CLK(clknet_1_0__leaf_wb_clk_i),
    .Q(\aaaa[8] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _237_ (.D(net90),
    .CLK(clknet_1_0__leaf_wb_clk_i),
    .Q(\aaaa[9] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _238_ (.D(net76),
    .CLK(clknet_1_1__leaf_wb_clk_i),
    .Q(\aaaa[10] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _239_ (.D(net77),
    .CLK(clknet_1_1__leaf_wb_clk_i),
    .Q(\aaaa[11] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _240_ (.D(net78),
    .CLK(clknet_1_1__leaf_wb_clk_i),
    .Q(\aaaa[12] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _241_ (.D(net79),
    .CLK(clknet_1_1__leaf_wb_clk_i),
    .Q(\aaaa[13] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _242_ (.D(net80),
    .CLK(clknet_1_1__leaf_wb_clk_i),
    .Q(\aaaa[14] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _243_ (.D(net81),
    .CLK(clknet_1_1__leaf_wb_clk_i),
    .Q(\aaaa[15] ));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 _252_ (.I(net84),
    .Z(net92));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _253_ (.I(net85),
    .Z(net93));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _254_ (.I(net86),
    .Z(net94));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _255_ (.I(net87),
    .Z(net95));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _256_ (.I(net88),
    .Z(net96));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _257_ (.I(net89),
    .Z(net97));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _258_ (.I(net90),
    .Z(net98));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _259_ (.I(net76),
    .Z(net99));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _260_ (.I(net77),
    .Z(net100));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _261_ (.I(net91),
    .Z(net101));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _262_ (.I(net66),
    .Z(net102));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _263_ (.I(net67),
    .Z(net103));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _264_ (.I(net68),
    .Z(net104));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _265_ (.I(net69),
    .Z(net105));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _266_ (.I(net70),
    .Z(net106));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _267_ (.I(net71),
    .Z(net107));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _268_ (.I(net72),
    .Z(net108));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _269_ (.I(net73),
    .Z(net109));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_0_wb_clk_i (.I(wb_clk_i),
    .Z(clknet_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_1_0__f_wb_clk_i (.I(clknet_0_wb_clk_i),
    .Z(clknet_1_0__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_1_1__f_wb_clk_i (.I(clknet_0_wb_clk_i),
    .Z(clknet_1_1__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 input1 (.I(Q0[0]),
    .Z(net1));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 input10 (.I(Q1[1]),
    .Z(net10));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 input11 (.I(Q1[2]),
    .Z(net11));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 input12 (.I(Q1[3]),
    .Z(net12));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 input13 (.I(Q1[4]),
    .Z(net13));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 input14 (.I(Q1[5]),
    .Z(net14));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input15 (.I(Q1[6]),
    .Z(net15));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input16 (.I(Q1[7]),
    .Z(net16));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 input17 (.I(Q2[0]),
    .Z(net17));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 input18 (.I(Q2[1]),
    .Z(net18));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 input19 (.I(Q2[2]),
    .Z(net19));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 input2 (.I(Q0[1]),
    .Z(net2));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 input20 (.I(Q2[3]),
    .Z(net20));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 input21 (.I(Q2[4]),
    .Z(net21));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input22 (.I(Q2[5]),
    .Z(net22));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 input23 (.I(Q2[6]),
    .Z(net23));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input24 (.I(Q2[7]),
    .Z(net24));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input25 (.I(Q3[0]),
    .Z(net25));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input26 (.I(Q3[1]),
    .Z(net26));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input27 (.I(Q3[2]),
    .Z(net27));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input28 (.I(Q3[3]),
    .Z(net28));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input29 (.I(Q3[4]),
    .Z(net29));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 input3 (.I(Q0[2]),
    .Z(net3));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input30 (.I(Q3[5]),
    .Z(net30));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input31 (.I(Q3[6]),
    .Z(net31));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input32 (.I(Q3[7]),
    .Z(net32));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input33 (.I(Q4[0]),
    .Z(net33));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input34 (.I(Q4[1]),
    .Z(net34));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input35 (.I(Q4[2]),
    .Z(net35));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input36 (.I(Q4[3]),
    .Z(net36));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input37 (.I(Q4[4]),
    .Z(net37));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input38 (.I(Q4[5]),
    .Z(net38));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 input39 (.I(Q4[6]),
    .Z(net39));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 input4 (.I(Q0[3]),
    .Z(net4));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 input40 (.I(Q4[7]),
    .Z(net40));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 input41 (.I(Q5[0]),
    .Z(net41));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 input42 (.I(Q5[1]),
    .Z(net42));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 input43 (.I(Q5[2]),
    .Z(net43));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 input44 (.I(Q5[3]),
    .Z(net44));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 input45 (.I(Q5[4]),
    .Z(net45));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 input46 (.I(Q5[5]),
    .Z(net46));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 input47 (.I(Q5[6]),
    .Z(net47));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 input48 (.I(Q5[7]),
    .Z(net48));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 input49 (.I(Q6[0]),
    .Z(net49));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 input5 (.I(Q0[4]),
    .Z(net5));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 input50 (.I(Q6[1]),
    .Z(net50));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 input51 (.I(Q6[2]),
    .Z(net51));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 input52 (.I(Q6[3]),
    .Z(net52));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 input53 (.I(Q6[4]),
    .Z(net53));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 input54 (.I(Q6[5]),
    .Z(net54));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 input55 (.I(Q6[6]),
    .Z(net55));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 input56 (.I(Q6[7]),
    .Z(net56));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 input57 (.I(Q7[0]),
    .Z(net57));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 input58 (.I(Q7[1]),
    .Z(net58));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 input59 (.I(Q7[2]),
    .Z(net59));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 input6 (.I(Q0[5]),
    .Z(net6));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 input60 (.I(Q7[3]),
    .Z(net60));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 input61 (.I(Q7[4]),
    .Z(net61));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 input62 (.I(Q7[5]),
    .Z(net62));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 input63 (.I(Q7[6]),
    .Z(net63));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 input64 (.I(Q7[7]),
    .Z(net64));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 input65 (.I(WEb_raw),
    .Z(net65));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 input66 (.I(bus_in[0]),
    .Z(net66));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 input67 (.I(bus_in[1]),
    .Z(net67));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 input68 (.I(bus_in[2]),
    .Z(net68));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 input69 (.I(bus_in[3]),
    .Z(net69));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 input7 (.I(Q0[6]),
    .Z(net7));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 input70 (.I(bus_in[4]),
    .Z(net70));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 input71 (.I(bus_in[5]),
    .Z(net71));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 input72 (.I(bus_in[6]),
    .Z(net72));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 input73 (.I(bus_in[7]),
    .Z(net73));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 input74 (.I(ram_enabled),
    .Z(net74));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 input75 (.I(requested_addr[0]),
    .Z(net75));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input76 (.I(requested_addr[10]),
    .Z(net76));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input77 (.I(requested_addr[11]),
    .Z(net77));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input78 (.I(requested_addr[12]),
    .Z(net78));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input79 (.I(requested_addr[13]),
    .Z(net79));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input8 (.I(Q0[7]),
    .Z(net8));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input80 (.I(requested_addr[14]),
    .Z(net80));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input81 (.I(requested_addr[15]),
    .Z(net81));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 input82 (.I(requested_addr[1]),
    .Z(net82));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 input83 (.I(requested_addr[2]),
    .Z(net83));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input84 (.I(requested_addr[3]),
    .Z(net84));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input85 (.I(requested_addr[4]),
    .Z(net85));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input86 (.I(requested_addr[5]),
    .Z(net86));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input87 (.I(requested_addr[6]),
    .Z(net87));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input88 (.I(requested_addr[7]),
    .Z(net88));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input89 (.I(requested_addr[8]),
    .Z(net89));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 input9 (.I(Q1[0]),
    .Z(net9));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input90 (.I(requested_addr[9]),
    .Z(net90));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 input91 (.I(rst),
    .Z(net91));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output100 (.I(net100),
    .Z(A_all[8]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output101 (.I(net101),
    .Z(CEN_all));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output102 (.I(net102),
    .Z(D_all[0]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output103 (.I(net103),
    .Z(D_all[1]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output104 (.I(net104),
    .Z(D_all[2]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output105 (.I(net105),
    .Z(D_all[3]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output106 (.I(net106),
    .Z(D_all[4]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output107 (.I(net107),
    .Z(D_all[5]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output108 (.I(net108),
    .Z(D_all[6]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output109 (.I(net109),
    .Z(D_all[7]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output110 (.I(net110),
    .Z(GWEN_0));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output111 (.I(net111),
    .Z(GWEN_1));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output112 (.I(net112),
    .Z(GWEN_2));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output113 (.I(net113),
    .Z(GWEN_3));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output114 (.I(net114),
    .Z(GWEN_4));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output115 (.I(net115),
    .Z(GWEN_5));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output116 (.I(net116),
    .Z(GWEN_6));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output117 (.I(net117),
    .Z(GWEN_7));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output118 (.I(net118),
    .Z(bus_out[0]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output119 (.I(net119),
    .Z(bus_out[1]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output120 (.I(net120),
    .Z(bus_out[2]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output121 (.I(net121),
    .Z(bus_out[3]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output122 (.I(net122),
    .Z(bus_out[4]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output123 (.I(net123),
    .Z(bus_out[5]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output124 (.I(net124),
    .Z(bus_out[6]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output125 (.I(net125),
    .Z(bus_out[7]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output92 (.I(net92),
    .Z(A_all[0]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output93 (.I(net93),
    .Z(A_all[1]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output94 (.I(net94),
    .Z(A_all[2]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output95 (.I(net95),
    .Z(A_all[3]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output96 (.I(net96),
    .Z(A_all[4]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output97 (.I(net97),
    .Z(A_all[5]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output98 (.I(net98),
    .Z(A_all[6]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output99 (.I(net99),
    .Z(A_all[7]));
 gf180mcu_fd_sc_mcu7t5v0__tiel ram_controller_126 (.ZN(net126));
 gf180mcu_fd_sc_mcu7t5v0__tiel ram_controller_127 (.ZN(net127));
 gf180mcu_fd_sc_mcu7t5v0__tiel ram_controller_128 (.ZN(net128));
 gf180mcu_fd_sc_mcu7t5v0__tiel ram_controller_129 (.ZN(net129));
 gf180mcu_fd_sc_mcu7t5v0__tiel ram_controller_130 (.ZN(net130));
 gf180mcu_fd_sc_mcu7t5v0__tiel ram_controller_131 (.ZN(net131));
 gf180mcu_fd_sc_mcu7t5v0__tiel ram_controller_132 (.ZN(net132));
 gf180mcu_fd_sc_mcu7t5v0__tiel ram_controller_133 (.ZN(net133));
 assign WEN_all[0] = net126;
 assign WEN_all[1] = net127;
 assign WEN_all[2] = net128;
 assign WEN_all[3] = net129;
 assign WEN_all[4] = net130;
 assign WEN_all[5] = net131;
 assign WEN_all[6] = net132;
 assign WEN_all[7] = net133;
endmodule

