VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO ram_controller
  CLASS BLOCK ;
  FOREIGN ram_controller ;
  ORIGIN 0.000 0.000 ;
  SIZE 1500.000 BY 300.000 ;
  PIN A_all[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 202.720 0.000 203.280 4.000 ;
    END
  END A_all[0]
  PIN A_all[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 220.640 0.000 221.200 4.000 ;
    END
  END A_all[1]
  PIN A_all[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 238.560 0.000 239.120 4.000 ;
    END
  END A_all[2]
  PIN A_all[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 256.480 0.000 257.040 4.000 ;
    END
  END A_all[3]
  PIN A_all[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 274.400 0.000 274.960 4.000 ;
    END
  END A_all[4]
  PIN A_all[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 292.320 0.000 292.880 4.000 ;
    END
  END A_all[5]
  PIN A_all[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 310.240 0.000 310.800 4.000 ;
    END
  END A_all[6]
  PIN A_all[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 328.160 0.000 328.720 4.000 ;
    END
  END A_all[7]
  PIN A_all[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 346.080 0.000 346.640 4.000 ;
    END
  END A_all[8]
  PIN CEN_all
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 41.440 0.000 42.000 4.000 ;
    END
  END CEN_all
  PIN D_all[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 364.000 0.000 364.560 4.000 ;
    END
  END D_all[0]
  PIN D_all[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 381.920 0.000 382.480 4.000 ;
    END
  END D_all[1]
  PIN D_all[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 399.840 0.000 400.400 4.000 ;
    END
  END D_all[2]
  PIN D_all[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 417.760 0.000 418.320 4.000 ;
    END
  END D_all[3]
  PIN D_all[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 435.680 0.000 436.240 4.000 ;
    END
  END D_all[4]
  PIN D_all[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 453.600 0.000 454.160 4.000 ;
    END
  END D_all[5]
  PIN D_all[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 471.520 0.000 472.080 4.000 ;
    END
  END D_all[6]
  PIN D_all[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 489.440 0.000 490.000 4.000 ;
    END
  END D_all[7]
  PIN GWEN_0
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 507.360 0.000 507.920 4.000 ;
    END
  END GWEN_0
  PIN GWEN_1
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 525.280 0.000 525.840 4.000 ;
    END
  END GWEN_1
  PIN GWEN_2
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 543.200 0.000 543.760 4.000 ;
    END
  END GWEN_2
  PIN GWEN_3
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 561.120 0.000 561.680 4.000 ;
    END
  END GWEN_3
  PIN GWEN_4
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 579.040 0.000 579.600 4.000 ;
    END
  END GWEN_4
  PIN GWEN_5
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 596.960 0.000 597.520 4.000 ;
    END
  END GWEN_5
  PIN GWEN_6
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 1004.640 296.000 1005.200 300.000 ;
    END
  END GWEN_6
  PIN GWEN_7
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 1031.520 296.000 1032.080 300.000 ;
    END
  END GWEN_7
  PIN Q0[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 614.880 0.000 615.440 4.000 ;
    END
  END Q0[0]
  PIN Q0[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 632.800 0.000 633.360 4.000 ;
    END
  END Q0[1]
  PIN Q0[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 650.720 0.000 651.280 4.000 ;
    END
  END Q0[2]
  PIN Q0[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 668.640 0.000 669.200 4.000 ;
    END
  END Q0[3]
  PIN Q0[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 686.560 0.000 687.120 4.000 ;
    END
  END Q0[4]
  PIN Q0[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 704.480 0.000 705.040 4.000 ;
    END
  END Q0[5]
  PIN Q0[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 722.400 0.000 722.960 4.000 ;
    END
  END Q0[6]
  PIN Q0[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 740.320 0.000 740.880 4.000 ;
    END
  END Q0[7]
  PIN Q1[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 758.240 0.000 758.800 4.000 ;
    END
  END Q1[0]
  PIN Q1[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 776.160 0.000 776.720 4.000 ;
    END
  END Q1[1]
  PIN Q1[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 794.080 0.000 794.640 4.000 ;
    END
  END Q1[2]
  PIN Q1[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 812.000 0.000 812.560 4.000 ;
    END
  END Q1[3]
  PIN Q1[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 829.920 0.000 830.480 4.000 ;
    END
  END Q1[4]
  PIN Q1[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 847.840 0.000 848.400 4.000 ;
    END
  END Q1[5]
  PIN Q1[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 865.760 0.000 866.320 4.000 ;
    END
  END Q1[6]
  PIN Q1[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 883.680 0.000 884.240 4.000 ;
    END
  END Q1[7]
  PIN Q2[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 901.600 0.000 902.160 4.000 ;
    END
  END Q2[0]
  PIN Q2[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 919.520 0.000 920.080 4.000 ;
    END
  END Q2[1]
  PIN Q2[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 937.440 0.000 938.000 4.000 ;
    END
  END Q2[2]
  PIN Q2[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 955.360 0.000 955.920 4.000 ;
    END
  END Q2[3]
  PIN Q2[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 973.280 0.000 973.840 4.000 ;
    END
  END Q2[4]
  PIN Q2[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 991.200 0.000 991.760 4.000 ;
    END
  END Q2[5]
  PIN Q2[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 1009.120 0.000 1009.680 4.000 ;
    END
  END Q2[6]
  PIN Q2[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 1027.040 0.000 1027.600 4.000 ;
    END
  END Q2[7]
  PIN Q3[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 1044.960 0.000 1045.520 4.000 ;
    END
  END Q3[0]
  PIN Q3[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 1062.880 0.000 1063.440 4.000 ;
    END
  END Q3[1]
  PIN Q3[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 1080.800 0.000 1081.360 4.000 ;
    END
  END Q3[2]
  PIN Q3[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 1098.720 0.000 1099.280 4.000 ;
    END
  END Q3[3]
  PIN Q3[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 1116.640 0.000 1117.200 4.000 ;
    END
  END Q3[4]
  PIN Q3[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 1134.560 0.000 1135.120 4.000 ;
    END
  END Q3[5]
  PIN Q3[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 1152.480 0.000 1153.040 4.000 ;
    END
  END Q3[6]
  PIN Q3[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 1170.400 0.000 1170.960 4.000 ;
    END
  END Q3[7]
  PIN Q4[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 1188.320 0.000 1188.880 4.000 ;
    END
  END Q4[0]
  PIN Q4[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 1206.240 0.000 1206.800 4.000 ;
    END
  END Q4[1]
  PIN Q4[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 1224.160 0.000 1224.720 4.000 ;
    END
  END Q4[2]
  PIN Q4[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 1242.080 0.000 1242.640 4.000 ;
    END
  END Q4[3]
  PIN Q4[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 1260.000 0.000 1260.560 4.000 ;
    END
  END Q4[4]
  PIN Q4[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 1277.920 0.000 1278.480 4.000 ;
    END
  END Q4[5]
  PIN Q4[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 1295.840 0.000 1296.400 4.000 ;
    END
  END Q4[6]
  PIN Q4[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 1313.760 0.000 1314.320 4.000 ;
    END
  END Q4[7]
  PIN Q5[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 1331.680 0.000 1332.240 4.000 ;
    END
  END Q5[0]
  PIN Q5[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 1349.600 0.000 1350.160 4.000 ;
    END
  END Q5[1]
  PIN Q5[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 1367.520 0.000 1368.080 4.000 ;
    END
  END Q5[2]
  PIN Q5[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 1385.440 0.000 1386.000 4.000 ;
    END
  END Q5[3]
  PIN Q5[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 1403.360 0.000 1403.920 4.000 ;
    END
  END Q5[4]
  PIN Q5[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 1421.280 0.000 1421.840 4.000 ;
    END
  END Q5[5]
  PIN Q5[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 1439.200 0.000 1439.760 4.000 ;
    END
  END Q5[6]
  PIN Q5[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 1457.120 0.000 1457.680 4.000 ;
    END
  END Q5[7]
  PIN Q6[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 1058.400 296.000 1058.960 300.000 ;
    END
  END Q6[0]
  PIN Q6[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 1085.280 296.000 1085.840 300.000 ;
    END
  END Q6[1]
  PIN Q6[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 1112.160 296.000 1112.720 300.000 ;
    END
  END Q6[2]
  PIN Q6[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 1139.040 296.000 1139.600 300.000 ;
    END
  END Q6[3]
  PIN Q6[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 1165.920 296.000 1166.480 300.000 ;
    END
  END Q6[4]
  PIN Q6[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.726000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 1192.800 296.000 1193.360 300.000 ;
    END
  END Q6[5]
  PIN Q6[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.726000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 1219.680 296.000 1220.240 300.000 ;
    END
  END Q6[6]
  PIN Q6[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.726000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 1246.560 296.000 1247.120 300.000 ;
    END
  END Q6[7]
  PIN Q7[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.183000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 1273.440 296.000 1274.000 300.000 ;
    END
  END Q7[0]
  PIN Q7[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.183000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 1300.320 296.000 1300.880 300.000 ;
    END
  END Q7[1]
  PIN Q7[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.183000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 1327.200 296.000 1327.760 300.000 ;
    END
  END Q7[2]
  PIN Q7[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.183000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 1354.080 296.000 1354.640 300.000 ;
    END
  END Q7[3]
  PIN Q7[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.183000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 1380.960 296.000 1381.520 300.000 ;
    END
  END Q7[4]
  PIN Q7[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.183000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 1407.840 296.000 1408.400 300.000 ;
    END
  END Q7[5]
  PIN Q7[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 1434.720 296.000 1435.280 300.000 ;
    END
  END Q7[6]
  PIN Q7[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 1461.600 296.000 1462.160 300.000 ;
    END
  END Q7[7]
  PIN WEN_all[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal2 ;
        RECT 59.360 0.000 59.920 4.000 ;
    END
  END WEN_all[0]
  PIN WEN_all[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal2 ;
        RECT 77.280 0.000 77.840 4.000 ;
    END
  END WEN_all[1]
  PIN WEN_all[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal2 ;
        RECT 95.200 0.000 95.760 4.000 ;
    END
  END WEN_all[2]
  PIN WEN_all[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal2 ;
        RECT 113.120 0.000 113.680 4.000 ;
    END
  END WEN_all[3]
  PIN WEN_all[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal2 ;
        RECT 131.040 0.000 131.600 4.000 ;
    END
  END WEN_all[4]
  PIN WEN_all[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal2 ;
        RECT 148.960 0.000 149.520 4.000 ;
    END
  END WEN_all[5]
  PIN WEN_all[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal2 ;
        RECT 166.880 0.000 167.440 4.000 ;
    END
  END WEN_all[6]
  PIN WEN_all[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal2 ;
        RECT 184.800 0.000 185.360 4.000 ;
    END
  END WEN_all[7]
  PIN WEb_raw
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 90.720 296.000 91.280 300.000 ;
    END
  END WEb_raw
  PIN bus_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 117.600 296.000 118.160 300.000 ;
    END
  END bus_in[0]
  PIN bus_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.726000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 144.480 296.000 145.040 300.000 ;
    END
  END bus_in[1]
  PIN bus_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.726000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 171.360 296.000 171.920 300.000 ;
    END
  END bus_in[2]
  PIN bus_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.726000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 198.240 296.000 198.800 300.000 ;
    END
  END bus_in[3]
  PIN bus_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.726000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 225.120 296.000 225.680 300.000 ;
    END
  END bus_in[4]
  PIN bus_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.726000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 252.000 296.000 252.560 300.000 ;
    END
  END bus_in[5]
  PIN bus_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.726000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 278.880 296.000 279.440 300.000 ;
    END
  END bus_in[6]
  PIN bus_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.726000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 305.760 296.000 306.320 300.000 ;
    END
  END bus_in[7]
  PIN bus_out[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 332.640 296.000 333.200 300.000 ;
    END
  END bus_out[0]
  PIN bus_out[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 359.520 296.000 360.080 300.000 ;
    END
  END bus_out[1]
  PIN bus_out[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 386.400 296.000 386.960 300.000 ;
    END
  END bus_out[2]
  PIN bus_out[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 413.280 296.000 413.840 300.000 ;
    END
  END bus_out[3]
  PIN bus_out[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 440.160 296.000 440.720 300.000 ;
    END
  END bus_out[4]
  PIN bus_out[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 467.040 296.000 467.600 300.000 ;
    END
  END bus_out[5]
  PIN bus_out[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 493.920 296.000 494.480 300.000 ;
    END
  END bus_out[6]
  PIN bus_out[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 520.800 296.000 521.360 300.000 ;
    END
  END bus_out[7]
  PIN ram_enabled
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.726000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 547.680 296.000 548.240 300.000 ;
    END
  END ram_enabled
  PIN requested_addr[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.726000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 574.560 296.000 575.120 300.000 ;
    END
  END requested_addr[0]
  PIN requested_addr[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 843.360 296.000 843.920 300.000 ;
    END
  END requested_addr[10]
  PIN requested_addr[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 870.240 296.000 870.800 300.000 ;
    END
  END requested_addr[11]
  PIN requested_addr[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 897.120 296.000 897.680 300.000 ;
    END
  END requested_addr[12]
  PIN requested_addr[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 924.000 296.000 924.560 300.000 ;
    END
  END requested_addr[13]
  PIN requested_addr[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 950.880 296.000 951.440 300.000 ;
    END
  END requested_addr[14]
  PIN requested_addr[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 977.760 296.000 978.320 300.000 ;
    END
  END requested_addr[15]
  PIN requested_addr[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.726000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 601.440 296.000 602.000 300.000 ;
    END
  END requested_addr[1]
  PIN requested_addr[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 628.320 296.000 628.880 300.000 ;
    END
  END requested_addr[2]
  PIN requested_addr[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 655.200 296.000 655.760 300.000 ;
    END
  END requested_addr[3]
  PIN requested_addr[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 682.080 296.000 682.640 300.000 ;
    END
  END requested_addr[4]
  PIN requested_addr[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 708.960 296.000 709.520 300.000 ;
    END
  END requested_addr[5]
  PIN requested_addr[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 735.840 296.000 736.400 300.000 ;
    END
  END requested_addr[6]
  PIN requested_addr[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 762.720 296.000 763.280 300.000 ;
    END
  END requested_addr[7]
  PIN requested_addr[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 789.600 296.000 790.160 300.000 ;
    END
  END requested_addr[8]
  PIN requested_addr[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 816.480 296.000 817.040 300.000 ;
    END
  END requested_addr[9]
  PIN rst
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 63.840 296.000 64.400 300.000 ;
    END
  END rst
  PIN vdd
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Metal4 ;
        RECT 22.240 15.380 23.840 282.540 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 175.840 15.380 177.440 282.540 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 329.440 15.380 331.040 282.540 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 483.040 15.380 484.640 282.540 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 636.640 15.380 638.240 282.540 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 790.240 15.380 791.840 282.540 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 943.840 15.380 945.440 282.540 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1097.440 15.380 1099.040 282.540 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1251.040 15.380 1252.640 282.540 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1404.640 15.380 1406.240 282.540 ;
    END
  END vdd
  PIN vss
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Metal4 ;
        RECT 99.040 15.380 100.640 282.540 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 252.640 15.380 254.240 282.540 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 406.240 15.380 407.840 282.540 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 559.840 15.380 561.440 282.540 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 713.440 15.380 715.040 282.540 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 867.040 15.380 868.640 282.540 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1020.640 15.380 1022.240 282.540 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1174.240 15.380 1175.840 282.540 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1327.840 15.380 1329.440 282.540 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1481.440 15.380 1483.040 282.540 ;
    END
  END vss
  PIN wb_clk_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 4.738000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 36.960 296.000 37.520 300.000 ;
    END
  END wb_clk_i
  OBS
      LAYER Pwell ;
        RECT 6.290 280.480 1493.390 282.670 ;
      LAYER Nwell ;
        RECT 6.290 276.285 1493.390 280.480 ;
        RECT 6.290 276.160 679.105 276.285 ;
      LAYER Pwell ;
        RECT 6.290 272.640 1493.390 276.160 ;
      LAYER Nwell ;
        RECT 6.290 272.515 657.480 272.640 ;
        RECT 6.290 268.445 1493.390 272.515 ;
        RECT 6.290 268.320 955.745 268.445 ;
      LAYER Pwell ;
        RECT 6.290 264.800 1493.390 268.320 ;
      LAYER Nwell ;
        RECT 6.290 264.675 916.545 264.800 ;
        RECT 6.290 260.480 1493.390 264.675 ;
      LAYER Pwell ;
        RECT 6.290 256.960 1493.390 260.480 ;
      LAYER Nwell ;
        RECT 6.290 252.640 1493.390 256.960 ;
      LAYER Pwell ;
        RECT 6.290 249.120 1493.390 252.640 ;
      LAYER Nwell ;
        RECT 6.290 244.800 1493.390 249.120 ;
      LAYER Pwell ;
        RECT 6.290 241.280 1493.390 244.800 ;
      LAYER Nwell ;
        RECT 6.290 236.960 1493.390 241.280 ;
      LAYER Pwell ;
        RECT 6.290 233.440 1493.390 236.960 ;
      LAYER Nwell ;
        RECT 6.290 229.120 1493.390 233.440 ;
      LAYER Pwell ;
        RECT 6.290 225.600 1493.390 229.120 ;
      LAYER Nwell ;
        RECT 6.290 221.280 1493.390 225.600 ;
      LAYER Pwell ;
        RECT 6.290 217.760 1493.390 221.280 ;
      LAYER Nwell ;
        RECT 6.290 213.440 1493.390 217.760 ;
      LAYER Pwell ;
        RECT 6.290 209.920 1493.390 213.440 ;
      LAYER Nwell ;
        RECT 6.290 205.600 1493.390 209.920 ;
      LAYER Pwell ;
        RECT 6.290 202.080 1493.390 205.600 ;
      LAYER Nwell ;
        RECT 6.290 197.760 1493.390 202.080 ;
      LAYER Pwell ;
        RECT 6.290 194.240 1493.390 197.760 ;
      LAYER Nwell ;
        RECT 6.290 189.920 1493.390 194.240 ;
      LAYER Pwell ;
        RECT 6.290 186.400 1493.390 189.920 ;
      LAYER Nwell ;
        RECT 6.290 182.080 1493.390 186.400 ;
      LAYER Pwell ;
        RECT 6.290 178.560 1493.390 182.080 ;
      LAYER Nwell ;
        RECT 6.290 174.240 1493.390 178.560 ;
      LAYER Pwell ;
        RECT 6.290 170.720 1493.390 174.240 ;
      LAYER Nwell ;
        RECT 6.290 166.400 1493.390 170.720 ;
      LAYER Pwell ;
        RECT 6.290 162.880 1493.390 166.400 ;
      LAYER Nwell ;
        RECT 6.290 158.560 1493.390 162.880 ;
      LAYER Pwell ;
        RECT 6.290 155.040 1493.390 158.560 ;
      LAYER Nwell ;
        RECT 6.290 150.720 1493.390 155.040 ;
      LAYER Pwell ;
        RECT 6.290 147.200 1493.390 150.720 ;
      LAYER Nwell ;
        RECT 6.290 142.880 1493.390 147.200 ;
      LAYER Pwell ;
        RECT 6.290 139.360 1493.390 142.880 ;
      LAYER Nwell ;
        RECT 6.290 135.040 1493.390 139.360 ;
      LAYER Pwell ;
        RECT 6.290 131.520 1493.390 135.040 ;
      LAYER Nwell ;
        RECT 6.290 127.200 1493.390 131.520 ;
      LAYER Pwell ;
        RECT 6.290 123.680 1493.390 127.200 ;
      LAYER Nwell ;
        RECT 6.290 119.360 1493.390 123.680 ;
      LAYER Pwell ;
        RECT 6.290 115.840 1493.390 119.360 ;
      LAYER Nwell ;
        RECT 6.290 111.520 1493.390 115.840 ;
      LAYER Pwell ;
        RECT 6.290 108.000 1493.390 111.520 ;
      LAYER Nwell ;
        RECT 6.290 103.680 1493.390 108.000 ;
      LAYER Pwell ;
        RECT 6.290 100.160 1493.390 103.680 ;
      LAYER Nwell ;
        RECT 6.290 95.840 1493.390 100.160 ;
      LAYER Pwell ;
        RECT 6.290 92.320 1493.390 95.840 ;
      LAYER Nwell ;
        RECT 6.290 88.000 1493.390 92.320 ;
      LAYER Pwell ;
        RECT 6.290 84.480 1493.390 88.000 ;
      LAYER Nwell ;
        RECT 6.290 80.160 1493.390 84.480 ;
      LAYER Pwell ;
        RECT 6.290 76.640 1493.390 80.160 ;
      LAYER Nwell ;
        RECT 6.290 72.320 1493.390 76.640 ;
      LAYER Pwell ;
        RECT 6.290 68.800 1493.390 72.320 ;
      LAYER Nwell ;
        RECT 6.290 64.480 1493.390 68.800 ;
      LAYER Pwell ;
        RECT 6.290 60.960 1493.390 64.480 ;
      LAYER Nwell ;
        RECT 6.290 56.640 1493.390 60.960 ;
      LAYER Pwell ;
        RECT 6.290 53.120 1493.390 56.640 ;
      LAYER Nwell ;
        RECT 6.290 48.800 1493.390 53.120 ;
      LAYER Pwell ;
        RECT 6.290 45.280 1493.390 48.800 ;
      LAYER Nwell ;
        RECT 6.290 45.155 963.025 45.280 ;
        RECT 6.290 40.960 1493.390 45.155 ;
      LAYER Pwell ;
        RECT 6.290 37.440 1493.390 40.960 ;
      LAYER Nwell ;
        RECT 6.290 37.315 926.625 37.440 ;
        RECT 6.290 33.120 1493.390 37.315 ;
      LAYER Pwell ;
        RECT 6.290 29.600 1493.390 33.120 ;
      LAYER Nwell ;
        RECT 6.290 29.475 917.105 29.600 ;
        RECT 6.290 25.405 1493.390 29.475 ;
        RECT 6.290 25.280 912.065 25.405 ;
      LAYER Pwell ;
        RECT 6.290 21.760 1493.390 25.280 ;
      LAYER Nwell ;
        RECT 6.290 21.635 917.105 21.760 ;
        RECT 6.290 17.565 1493.390 21.635 ;
        RECT 6.290 17.440 961.905 17.565 ;
      LAYER Pwell ;
        RECT 6.290 15.250 1493.390 17.440 ;
      LAYER Metal1 ;
        RECT 6.720 15.380 1492.960 285.450 ;
      LAYER Metal2 ;
        RECT 22.380 295.700 36.660 296.000 ;
        RECT 37.820 295.700 63.540 296.000 ;
        RECT 64.700 295.700 90.420 296.000 ;
        RECT 91.580 295.700 117.300 296.000 ;
        RECT 118.460 295.700 144.180 296.000 ;
        RECT 145.340 295.700 171.060 296.000 ;
        RECT 172.220 295.700 197.940 296.000 ;
        RECT 199.100 295.700 224.820 296.000 ;
        RECT 225.980 295.700 251.700 296.000 ;
        RECT 252.860 295.700 278.580 296.000 ;
        RECT 279.740 295.700 305.460 296.000 ;
        RECT 306.620 295.700 332.340 296.000 ;
        RECT 333.500 295.700 359.220 296.000 ;
        RECT 360.380 295.700 386.100 296.000 ;
        RECT 387.260 295.700 412.980 296.000 ;
        RECT 414.140 295.700 439.860 296.000 ;
        RECT 441.020 295.700 466.740 296.000 ;
        RECT 467.900 295.700 493.620 296.000 ;
        RECT 494.780 295.700 520.500 296.000 ;
        RECT 521.660 295.700 547.380 296.000 ;
        RECT 548.540 295.700 574.260 296.000 ;
        RECT 575.420 295.700 601.140 296.000 ;
        RECT 602.300 295.700 628.020 296.000 ;
        RECT 629.180 295.700 654.900 296.000 ;
        RECT 656.060 295.700 681.780 296.000 ;
        RECT 682.940 295.700 708.660 296.000 ;
        RECT 709.820 295.700 735.540 296.000 ;
        RECT 736.700 295.700 762.420 296.000 ;
        RECT 763.580 295.700 789.300 296.000 ;
        RECT 790.460 295.700 816.180 296.000 ;
        RECT 817.340 295.700 843.060 296.000 ;
        RECT 844.220 295.700 869.940 296.000 ;
        RECT 871.100 295.700 896.820 296.000 ;
        RECT 897.980 295.700 923.700 296.000 ;
        RECT 924.860 295.700 950.580 296.000 ;
        RECT 951.740 295.700 977.460 296.000 ;
        RECT 978.620 295.700 1004.340 296.000 ;
        RECT 1005.500 295.700 1031.220 296.000 ;
        RECT 1032.380 295.700 1058.100 296.000 ;
        RECT 1059.260 295.700 1084.980 296.000 ;
        RECT 1086.140 295.700 1111.860 296.000 ;
        RECT 1113.020 295.700 1138.740 296.000 ;
        RECT 1139.900 295.700 1165.620 296.000 ;
        RECT 1166.780 295.700 1192.500 296.000 ;
        RECT 1193.660 295.700 1219.380 296.000 ;
        RECT 1220.540 295.700 1246.260 296.000 ;
        RECT 1247.420 295.700 1273.140 296.000 ;
        RECT 1274.300 295.700 1300.020 296.000 ;
        RECT 1301.180 295.700 1326.900 296.000 ;
        RECT 1328.060 295.700 1353.780 296.000 ;
        RECT 1354.940 295.700 1380.660 296.000 ;
        RECT 1381.820 295.700 1407.540 296.000 ;
        RECT 1408.700 295.700 1434.420 296.000 ;
        RECT 1435.580 295.700 1461.300 296.000 ;
        RECT 1462.460 295.700 1482.900 296.000 ;
        RECT 22.380 4.300 1482.900 295.700 ;
        RECT 22.380 3.500 41.140 4.300 ;
        RECT 42.300 3.500 59.060 4.300 ;
        RECT 60.220 3.500 76.980 4.300 ;
        RECT 78.140 3.500 94.900 4.300 ;
        RECT 96.060 3.500 112.820 4.300 ;
        RECT 113.980 3.500 130.740 4.300 ;
        RECT 131.900 3.500 148.660 4.300 ;
        RECT 149.820 3.500 166.580 4.300 ;
        RECT 167.740 3.500 184.500 4.300 ;
        RECT 185.660 3.500 202.420 4.300 ;
        RECT 203.580 3.500 220.340 4.300 ;
        RECT 221.500 3.500 238.260 4.300 ;
        RECT 239.420 3.500 256.180 4.300 ;
        RECT 257.340 3.500 274.100 4.300 ;
        RECT 275.260 3.500 292.020 4.300 ;
        RECT 293.180 3.500 309.940 4.300 ;
        RECT 311.100 3.500 327.860 4.300 ;
        RECT 329.020 3.500 345.780 4.300 ;
        RECT 346.940 3.500 363.700 4.300 ;
        RECT 364.860 3.500 381.620 4.300 ;
        RECT 382.780 3.500 399.540 4.300 ;
        RECT 400.700 3.500 417.460 4.300 ;
        RECT 418.620 3.500 435.380 4.300 ;
        RECT 436.540 3.500 453.300 4.300 ;
        RECT 454.460 3.500 471.220 4.300 ;
        RECT 472.380 3.500 489.140 4.300 ;
        RECT 490.300 3.500 507.060 4.300 ;
        RECT 508.220 3.500 524.980 4.300 ;
        RECT 526.140 3.500 542.900 4.300 ;
        RECT 544.060 3.500 560.820 4.300 ;
        RECT 561.980 3.500 578.740 4.300 ;
        RECT 579.900 3.500 596.660 4.300 ;
        RECT 597.820 3.500 614.580 4.300 ;
        RECT 615.740 3.500 632.500 4.300 ;
        RECT 633.660 3.500 650.420 4.300 ;
        RECT 651.580 3.500 668.340 4.300 ;
        RECT 669.500 3.500 686.260 4.300 ;
        RECT 687.420 3.500 704.180 4.300 ;
        RECT 705.340 3.500 722.100 4.300 ;
        RECT 723.260 3.500 740.020 4.300 ;
        RECT 741.180 3.500 757.940 4.300 ;
        RECT 759.100 3.500 775.860 4.300 ;
        RECT 777.020 3.500 793.780 4.300 ;
        RECT 794.940 3.500 811.700 4.300 ;
        RECT 812.860 3.500 829.620 4.300 ;
        RECT 830.780 3.500 847.540 4.300 ;
        RECT 848.700 3.500 865.460 4.300 ;
        RECT 866.620 3.500 883.380 4.300 ;
        RECT 884.540 3.500 901.300 4.300 ;
        RECT 902.460 3.500 919.220 4.300 ;
        RECT 920.380 3.500 937.140 4.300 ;
        RECT 938.300 3.500 955.060 4.300 ;
        RECT 956.220 3.500 972.980 4.300 ;
        RECT 974.140 3.500 990.900 4.300 ;
        RECT 992.060 3.500 1008.820 4.300 ;
        RECT 1009.980 3.500 1026.740 4.300 ;
        RECT 1027.900 3.500 1044.660 4.300 ;
        RECT 1045.820 3.500 1062.580 4.300 ;
        RECT 1063.740 3.500 1080.500 4.300 ;
        RECT 1081.660 3.500 1098.420 4.300 ;
        RECT 1099.580 3.500 1116.340 4.300 ;
        RECT 1117.500 3.500 1134.260 4.300 ;
        RECT 1135.420 3.500 1152.180 4.300 ;
        RECT 1153.340 3.500 1170.100 4.300 ;
        RECT 1171.260 3.500 1188.020 4.300 ;
        RECT 1189.180 3.500 1205.940 4.300 ;
        RECT 1207.100 3.500 1223.860 4.300 ;
        RECT 1225.020 3.500 1241.780 4.300 ;
        RECT 1242.940 3.500 1259.700 4.300 ;
        RECT 1260.860 3.500 1277.620 4.300 ;
        RECT 1278.780 3.500 1295.540 4.300 ;
        RECT 1296.700 3.500 1313.460 4.300 ;
        RECT 1314.620 3.500 1331.380 4.300 ;
        RECT 1332.540 3.500 1349.300 4.300 ;
        RECT 1350.460 3.500 1367.220 4.300 ;
        RECT 1368.380 3.500 1385.140 4.300 ;
        RECT 1386.300 3.500 1403.060 4.300 ;
        RECT 1404.220 3.500 1420.980 4.300 ;
        RECT 1422.140 3.500 1438.900 4.300 ;
        RECT 1440.060 3.500 1456.820 4.300 ;
        RECT 1457.980 3.500 1482.900 4.300 ;
      LAYER Metal3 ;
        RECT 22.330 5.180 1482.950 282.380 ;
      LAYER Metal4 ;
        RECT 1085.420 22.490 1097.140 52.550 ;
        RECT 1099.340 22.490 1104.180 52.550 ;
  END
END ram_controller
END LIBRARY

