VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO ram_controller
  CLASS BLOCK ;
  FOREIGN ram_controller ;
  ORIGIN 0.000 0.000 ;
  SIZE 1100.000 BY 250.000 ;
  PIN A_all[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 138.880 0.000 139.440 4.000 ;
    END
  END A_all[0]
  PIN A_all[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 152.320 0.000 152.880 4.000 ;
    END
  END A_all[1]
  PIN A_all[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 165.760 0.000 166.320 4.000 ;
    END
  END A_all[2]
  PIN A_all[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 179.200 0.000 179.760 4.000 ;
    END
  END A_all[3]
  PIN A_all[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 192.640 0.000 193.200 4.000 ;
    END
  END A_all[4]
  PIN A_all[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 206.080 0.000 206.640 4.000 ;
    END
  END A_all[5]
  PIN A_all[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 219.520 0.000 220.080 4.000 ;
    END
  END A_all[6]
  PIN A_all[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 232.960 0.000 233.520 4.000 ;
    END
  END A_all[7]
  PIN A_all[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 246.400 0.000 246.960 4.000 ;
    END
  END A_all[8]
  PIN CEN_all
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 17.920 0.000 18.480 4.000 ;
    END
  END CEN_all
  PIN D_all[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 259.840 0.000 260.400 4.000 ;
    END
  END D_all[0]
  PIN D_all[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 273.280 0.000 273.840 4.000 ;
    END
  END D_all[1]
  PIN D_all[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 286.720 0.000 287.280 4.000 ;
    END
  END D_all[2]
  PIN D_all[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 300.160 0.000 300.720 4.000 ;
    END
  END D_all[3]
  PIN D_all[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 313.600 0.000 314.160 4.000 ;
    END
  END D_all[4]
  PIN D_all[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 327.040 0.000 327.600 4.000 ;
    END
  END D_all[5]
  PIN D_all[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 340.480 0.000 341.040 4.000 ;
    END
  END D_all[6]
  PIN D_all[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 353.920 0.000 354.480 4.000 ;
    END
  END D_all[7]
  PIN GWEN_0
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 367.360 0.000 367.920 4.000 ;
    END
  END GWEN_0
  PIN GWEN_1
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 380.800 0.000 381.360 4.000 ;
    END
  END GWEN_1
  PIN GWEN_2
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 394.240 0.000 394.800 4.000 ;
    END
  END GWEN_2
  PIN GWEN_3
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 407.680 0.000 408.240 4.000 ;
    END
  END GWEN_3
  PIN GWEN_4
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 421.120 0.000 421.680 4.000 ;
    END
  END GWEN_4
  PIN GWEN_5
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 434.560 0.000 435.120 4.000 ;
    END
  END GWEN_5
  PIN GWEN_6
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 740.320 246.000 740.880 250.000 ;
    END
  END GWEN_6
  PIN GWEN_7
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 760.480 246.000 761.040 250.000 ;
    END
  END GWEN_7
  PIN Q0[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 448.000 0.000 448.560 4.000 ;
    END
  END Q0[0]
  PIN Q0[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 461.440 0.000 462.000 4.000 ;
    END
  END Q0[1]
  PIN Q0[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 474.880 0.000 475.440 4.000 ;
    END
  END Q0[2]
  PIN Q0[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 488.320 0.000 488.880 4.000 ;
    END
  END Q0[3]
  PIN Q0[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 501.760 0.000 502.320 4.000 ;
    END
  END Q0[4]
  PIN Q0[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 515.200 0.000 515.760 4.000 ;
    END
  END Q0[5]
  PIN Q0[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 528.640 0.000 529.200 4.000 ;
    END
  END Q0[6]
  PIN Q0[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 542.080 0.000 542.640 4.000 ;
    END
  END Q0[7]
  PIN Q1[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 555.520 0.000 556.080 4.000 ;
    END
  END Q1[0]
  PIN Q1[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 568.960 0.000 569.520 4.000 ;
    END
  END Q1[1]
  PIN Q1[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 582.400 0.000 582.960 4.000 ;
    END
  END Q1[2]
  PIN Q1[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 595.840 0.000 596.400 4.000 ;
    END
  END Q1[3]
  PIN Q1[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 609.280 0.000 609.840 4.000 ;
    END
  END Q1[4]
  PIN Q1[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 622.720 0.000 623.280 4.000 ;
    END
  END Q1[5]
  PIN Q1[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 636.160 0.000 636.720 4.000 ;
    END
  END Q1[6]
  PIN Q1[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 649.600 0.000 650.160 4.000 ;
    END
  END Q1[7]
  PIN Q2[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 663.040 0.000 663.600 4.000 ;
    END
  END Q2[0]
  PIN Q2[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 676.480 0.000 677.040 4.000 ;
    END
  END Q2[1]
  PIN Q2[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 689.920 0.000 690.480 4.000 ;
    END
  END Q2[2]
  PIN Q2[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 703.360 0.000 703.920 4.000 ;
    END
  END Q2[3]
  PIN Q2[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 716.800 0.000 717.360 4.000 ;
    END
  END Q2[4]
  PIN Q2[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 730.240 0.000 730.800 4.000 ;
    END
  END Q2[5]
  PIN Q2[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 743.680 0.000 744.240 4.000 ;
    END
  END Q2[6]
  PIN Q2[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 757.120 0.000 757.680 4.000 ;
    END
  END Q2[7]
  PIN Q3[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 770.560 0.000 771.120 4.000 ;
    END
  END Q3[0]
  PIN Q3[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 784.000 0.000 784.560 4.000 ;
    END
  END Q3[1]
  PIN Q3[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 797.440 0.000 798.000 4.000 ;
    END
  END Q3[2]
  PIN Q3[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 810.880 0.000 811.440 4.000 ;
    END
  END Q3[3]
  PIN Q3[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 824.320 0.000 824.880 4.000 ;
    END
  END Q3[4]
  PIN Q3[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 837.760 0.000 838.320 4.000 ;
    END
  END Q3[5]
  PIN Q3[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 851.200 0.000 851.760 4.000 ;
    END
  END Q3[6]
  PIN Q3[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 864.640 0.000 865.200 4.000 ;
    END
  END Q3[7]
  PIN Q4[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 878.080 0.000 878.640 4.000 ;
    END
  END Q4[0]
  PIN Q4[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 891.520 0.000 892.080 4.000 ;
    END
  END Q4[1]
  PIN Q4[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 904.960 0.000 905.520 4.000 ;
    END
  END Q4[2]
  PIN Q4[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 918.400 0.000 918.960 4.000 ;
    END
  END Q4[3]
  PIN Q4[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 931.840 0.000 932.400 4.000 ;
    END
  END Q4[4]
  PIN Q4[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 945.280 0.000 945.840 4.000 ;
    END
  END Q4[5]
  PIN Q4[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 958.720 0.000 959.280 4.000 ;
    END
  END Q4[6]
  PIN Q4[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 972.160 0.000 972.720 4.000 ;
    END
  END Q4[7]
  PIN Q5[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.726000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 985.600 0.000 986.160 4.000 ;
    END
  END Q5[0]
  PIN Q5[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 999.040 0.000 999.600 4.000 ;
    END
  END Q5[1]
  PIN Q5[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 1012.480 0.000 1013.040 4.000 ;
    END
  END Q5[2]
  PIN Q5[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.726000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 1025.920 0.000 1026.480 4.000 ;
    END
  END Q5[3]
  PIN Q5[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 1039.360 0.000 1039.920 4.000 ;
    END
  END Q5[4]
  PIN Q5[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 1052.800 0.000 1053.360 4.000 ;
    END
  END Q5[5]
  PIN Q5[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 1066.240 0.000 1066.800 4.000 ;
    END
  END Q5[6]
  PIN Q5[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 1079.680 0.000 1080.240 4.000 ;
    END
  END Q5[7]
  PIN Q6[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 780.640 246.000 781.200 250.000 ;
    END
  END Q6[0]
  PIN Q6[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 800.800 246.000 801.360 250.000 ;
    END
  END Q6[1]
  PIN Q6[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 820.960 246.000 821.520 250.000 ;
    END
  END Q6[2]
  PIN Q6[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 841.120 246.000 841.680 250.000 ;
    END
  END Q6[3]
  PIN Q6[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 861.280 246.000 861.840 250.000 ;
    END
  END Q6[4]
  PIN Q6[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 881.440 246.000 882.000 250.000 ;
    END
  END Q6[5]
  PIN Q6[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 901.600 246.000 902.160 250.000 ;
    END
  END Q6[6]
  PIN Q6[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 921.760 246.000 922.320 250.000 ;
    END
  END Q6[7]
  PIN Q7[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 941.920 246.000 942.480 250.000 ;
    END
  END Q7[0]
  PIN Q7[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 962.080 246.000 962.640 250.000 ;
    END
  END Q7[1]
  PIN Q7[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 982.240 246.000 982.800 250.000 ;
    END
  END Q7[2]
  PIN Q7[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 1002.400 246.000 1002.960 250.000 ;
    END
  END Q7[3]
  PIN Q7[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 1022.560 246.000 1023.120 250.000 ;
    END
  END Q7[4]
  PIN Q7[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 1042.720 246.000 1043.280 250.000 ;
    END
  END Q7[5]
  PIN Q7[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.183000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 1062.880 246.000 1063.440 250.000 ;
    END
  END Q7[6]
  PIN Q7[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.183000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 1083.040 246.000 1083.600 250.000 ;
    END
  END Q7[7]
  PIN WEN_all[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal2 ;
        RECT 31.360 0.000 31.920 4.000 ;
    END
  END WEN_all[0]
  PIN WEN_all[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal2 ;
        RECT 44.800 0.000 45.360 4.000 ;
    END
  END WEN_all[1]
  PIN WEN_all[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal2 ;
        RECT 58.240 0.000 58.800 4.000 ;
    END
  END WEN_all[2]
  PIN WEN_all[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal2 ;
        RECT 71.680 0.000 72.240 4.000 ;
    END
  END WEN_all[3]
  PIN WEN_all[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal2 ;
        RECT 85.120 0.000 85.680 4.000 ;
    END
  END WEN_all[4]
  PIN WEN_all[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal2 ;
        RECT 98.560 0.000 99.120 4.000 ;
    END
  END WEN_all[5]
  PIN WEN_all[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal2 ;
        RECT 112.000 0.000 112.560 4.000 ;
    END
  END WEN_all[6]
  PIN WEN_all[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal2 ;
        RECT 125.440 0.000 126.000 4.000 ;
    END
  END WEN_all[7]
  PIN WEb_ram
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.183000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 54.880 246.000 55.440 250.000 ;
    END
  END WEb_ram
  PIN bus_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.726000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 75.040 246.000 75.600 250.000 ;
    END
  END bus_in[0]
  PIN bus_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.726000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 95.200 246.000 95.760 250.000 ;
    END
  END bus_in[1]
  PIN bus_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.726000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 115.360 246.000 115.920 250.000 ;
    END
  END bus_in[2]
  PIN bus_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.726000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 135.520 246.000 136.080 250.000 ;
    END
  END bus_in[3]
  PIN bus_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.726000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 155.680 246.000 156.240 250.000 ;
    END
  END bus_in[4]
  PIN bus_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.726000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 175.840 246.000 176.400 250.000 ;
    END
  END bus_in[5]
  PIN bus_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.726000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 196.000 246.000 196.560 250.000 ;
    END
  END bus_in[6]
  PIN bus_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.726000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 216.160 246.000 216.720 250.000 ;
    END
  END bus_in[7]
  PIN bus_out[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 236.320 246.000 236.880 250.000 ;
    END
  END bus_out[0]
  PIN bus_out[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 256.480 246.000 257.040 250.000 ;
    END
  END bus_out[1]
  PIN bus_out[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 276.640 246.000 277.200 250.000 ;
    END
  END bus_out[2]
  PIN bus_out[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 296.800 246.000 297.360 250.000 ;
    END
  END bus_out[3]
  PIN bus_out[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 316.960 246.000 317.520 250.000 ;
    END
  END bus_out[4]
  PIN bus_out[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 337.120 246.000 337.680 250.000 ;
    END
  END bus_out[5]
  PIN bus_out[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 357.280 246.000 357.840 250.000 ;
    END
  END bus_out[6]
  PIN bus_out[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 377.440 246.000 378.000 250.000 ;
    END
  END bus_out[7]
  PIN ram_enabled
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 397.600 246.000 398.160 250.000 ;
    END
  END ram_enabled
  PIN requested_addr[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 417.760 246.000 418.320 250.000 ;
    END
  END requested_addr[0]
  PIN requested_addr[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 619.360 246.000 619.920 250.000 ;
    END
  END requested_addr[10]
  PIN requested_addr[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 639.520 246.000 640.080 250.000 ;
    END
  END requested_addr[11]
  PIN requested_addr[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 659.680 246.000 660.240 250.000 ;
    END
  END requested_addr[12]
  PIN requested_addr[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 679.840 246.000 680.400 250.000 ;
    END
  END requested_addr[13]
  PIN requested_addr[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 700.000 246.000 700.560 250.000 ;
    END
  END requested_addr[14]
  PIN requested_addr[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 720.160 246.000 720.720 250.000 ;
    END
  END requested_addr[15]
  PIN requested_addr[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 437.920 246.000 438.480 250.000 ;
    END
  END requested_addr[1]
  PIN requested_addr[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 458.080 246.000 458.640 250.000 ;
    END
  END requested_addr[2]
  PIN requested_addr[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 478.240 246.000 478.800 250.000 ;
    END
  END requested_addr[3]
  PIN requested_addr[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 498.400 246.000 498.960 250.000 ;
    END
  END requested_addr[4]
  PIN requested_addr[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 518.560 246.000 519.120 250.000 ;
    END
  END requested_addr[5]
  PIN requested_addr[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 538.720 246.000 539.280 250.000 ;
    END
  END requested_addr[6]
  PIN requested_addr[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 558.880 246.000 559.440 250.000 ;
    END
  END requested_addr[7]
  PIN requested_addr[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 579.040 246.000 579.600 250.000 ;
    END
  END requested_addr[8]
  PIN requested_addr[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 599.200 246.000 599.760 250.000 ;
    END
  END requested_addr[9]
  PIN rst
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 34.720 246.000 35.280 250.000 ;
    END
  END rst
  PIN vdd
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Metal4 ;
        RECT 22.240 15.380 23.840 231.580 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 175.840 15.380 177.440 231.580 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 329.440 15.380 331.040 231.580 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 483.040 15.380 484.640 231.580 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 636.640 15.380 638.240 231.580 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 790.240 15.380 791.840 231.580 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 943.840 15.380 945.440 231.580 ;
    END
  END vdd
  PIN vss
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Metal4 ;
        RECT 99.040 15.380 100.640 231.580 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 252.640 15.380 254.240 231.580 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 406.240 15.380 407.840 231.580 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 559.840 15.380 561.440 231.580 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 713.440 15.380 715.040 231.580 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 867.040 15.380 868.640 231.580 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1020.640 15.380 1022.240 231.580 ;
    END
  END vss
  PIN wb_clk_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 4.738000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 14.560 246.000 15.120 250.000 ;
    END
  END wb_clk_i
  OBS
      LAYER Nwell ;
        RECT 6.290 229.120 1093.550 231.710 ;
      LAYER Pwell ;
        RECT 6.290 225.600 1093.550 229.120 ;
      LAYER Nwell ;
        RECT 6.290 221.405 1093.550 225.600 ;
        RECT 6.290 221.280 663.425 221.405 ;
      LAYER Pwell ;
        RECT 6.290 217.760 1093.550 221.280 ;
      LAYER Nwell ;
        RECT 6.290 217.635 697.240 217.760 ;
        RECT 6.290 213.440 1093.550 217.635 ;
      LAYER Pwell ;
        RECT 6.290 209.920 1093.550 213.440 ;
      LAYER Nwell ;
        RECT 6.290 205.600 1093.550 209.920 ;
      LAYER Pwell ;
        RECT 6.290 202.080 1093.550 205.600 ;
      LAYER Nwell ;
        RECT 6.290 197.760 1093.550 202.080 ;
      LAYER Pwell ;
        RECT 6.290 194.240 1093.550 197.760 ;
      LAYER Nwell ;
        RECT 6.290 189.920 1093.550 194.240 ;
      LAYER Pwell ;
        RECT 6.290 186.400 1093.550 189.920 ;
      LAYER Nwell ;
        RECT 6.290 182.080 1093.550 186.400 ;
      LAYER Pwell ;
        RECT 6.290 178.560 1093.550 182.080 ;
      LAYER Nwell ;
        RECT 6.290 174.240 1093.550 178.560 ;
      LAYER Pwell ;
        RECT 6.290 170.720 1093.550 174.240 ;
      LAYER Nwell ;
        RECT 6.290 166.400 1093.550 170.720 ;
      LAYER Pwell ;
        RECT 6.290 162.880 1093.550 166.400 ;
      LAYER Nwell ;
        RECT 6.290 158.560 1093.550 162.880 ;
      LAYER Pwell ;
        RECT 6.290 155.040 1093.550 158.560 ;
      LAYER Nwell ;
        RECT 6.290 154.915 539.880 155.040 ;
        RECT 6.290 150.845 1093.550 154.915 ;
        RECT 6.290 150.720 476.040 150.845 ;
      LAYER Pwell ;
        RECT 6.290 147.200 1093.550 150.720 ;
      LAYER Nwell ;
        RECT 6.290 147.075 499.000 147.200 ;
        RECT 6.290 142.880 1093.550 147.075 ;
      LAYER Pwell ;
        RECT 6.290 139.360 1093.550 142.880 ;
      LAYER Nwell ;
        RECT 6.290 135.040 1093.550 139.360 ;
      LAYER Pwell ;
        RECT 6.290 131.520 1093.550 135.040 ;
      LAYER Nwell ;
        RECT 6.290 127.200 1093.550 131.520 ;
      LAYER Pwell ;
        RECT 6.290 123.680 1093.550 127.200 ;
      LAYER Nwell ;
        RECT 6.290 119.360 1093.550 123.680 ;
      LAYER Pwell ;
        RECT 6.290 115.840 1093.550 119.360 ;
      LAYER Nwell ;
        RECT 6.290 111.520 1093.550 115.840 ;
      LAYER Pwell ;
        RECT 6.290 108.000 1093.550 111.520 ;
      LAYER Nwell ;
        RECT 6.290 103.680 1093.550 108.000 ;
      LAYER Pwell ;
        RECT 6.290 100.160 1093.550 103.680 ;
      LAYER Nwell ;
        RECT 6.290 95.840 1093.550 100.160 ;
      LAYER Pwell ;
        RECT 6.290 92.320 1093.550 95.840 ;
      LAYER Nwell ;
        RECT 6.290 88.000 1093.550 92.320 ;
      LAYER Pwell ;
        RECT 6.290 84.480 1093.550 88.000 ;
      LAYER Nwell ;
        RECT 6.290 80.160 1093.550 84.480 ;
      LAYER Pwell ;
        RECT 6.290 76.640 1093.550 80.160 ;
      LAYER Nwell ;
        RECT 6.290 72.320 1093.550 76.640 ;
      LAYER Pwell ;
        RECT 6.290 68.800 1093.550 72.320 ;
      LAYER Nwell ;
        RECT 6.290 64.480 1093.550 68.800 ;
      LAYER Pwell ;
        RECT 6.290 60.960 1093.550 64.480 ;
      LAYER Nwell ;
        RECT 6.290 56.640 1093.550 60.960 ;
      LAYER Pwell ;
        RECT 6.290 53.120 1093.550 56.640 ;
      LAYER Nwell ;
        RECT 6.290 52.995 781.350 53.120 ;
        RECT 6.290 48.800 1093.550 52.995 ;
      LAYER Pwell ;
        RECT 6.290 45.280 1093.550 48.800 ;
      LAYER Nwell ;
        RECT 6.290 45.155 676.305 45.280 ;
        RECT 6.290 41.085 1093.550 45.155 ;
        RECT 6.290 40.960 663.985 41.085 ;
      LAYER Pwell ;
        RECT 6.290 37.440 1093.550 40.960 ;
      LAYER Nwell ;
        RECT 6.290 37.315 657.265 37.440 ;
        RECT 6.290 33.245 1093.550 37.315 ;
        RECT 6.290 33.120 663.985 33.245 ;
      LAYER Pwell ;
        RECT 6.290 29.600 1093.550 33.120 ;
      LAYER Nwell ;
        RECT 6.290 29.475 680.785 29.600 ;
        RECT 6.290 25.280 1093.550 29.475 ;
      LAYER Pwell ;
        RECT 6.290 21.760 1093.550 25.280 ;
      LAYER Nwell ;
        RECT 6.290 21.635 758.070 21.760 ;
        RECT 6.290 17.440 1093.550 21.635 ;
      LAYER Pwell ;
        RECT 6.290 15.250 1093.550 17.440 ;
      LAYER Metal1 ;
        RECT 6.720 15.380 1093.120 232.250 ;
      LAYER Metal2 ;
        RECT 15.420 245.700 34.420 246.000 ;
        RECT 35.580 245.700 54.580 246.000 ;
        RECT 55.740 245.700 74.740 246.000 ;
        RECT 75.900 245.700 94.900 246.000 ;
        RECT 96.060 245.700 115.060 246.000 ;
        RECT 116.220 245.700 135.220 246.000 ;
        RECT 136.380 245.700 155.380 246.000 ;
        RECT 156.540 245.700 175.540 246.000 ;
        RECT 176.700 245.700 195.700 246.000 ;
        RECT 196.860 245.700 215.860 246.000 ;
        RECT 217.020 245.700 236.020 246.000 ;
        RECT 237.180 245.700 256.180 246.000 ;
        RECT 257.340 245.700 276.340 246.000 ;
        RECT 277.500 245.700 296.500 246.000 ;
        RECT 297.660 245.700 316.660 246.000 ;
        RECT 317.820 245.700 336.820 246.000 ;
        RECT 337.980 245.700 356.980 246.000 ;
        RECT 358.140 245.700 377.140 246.000 ;
        RECT 378.300 245.700 397.300 246.000 ;
        RECT 398.460 245.700 417.460 246.000 ;
        RECT 418.620 245.700 437.620 246.000 ;
        RECT 438.780 245.700 457.780 246.000 ;
        RECT 458.940 245.700 477.940 246.000 ;
        RECT 479.100 245.700 498.100 246.000 ;
        RECT 499.260 245.700 518.260 246.000 ;
        RECT 519.420 245.700 538.420 246.000 ;
        RECT 539.580 245.700 558.580 246.000 ;
        RECT 559.740 245.700 578.740 246.000 ;
        RECT 579.900 245.700 598.900 246.000 ;
        RECT 600.060 245.700 619.060 246.000 ;
        RECT 620.220 245.700 639.220 246.000 ;
        RECT 640.380 245.700 659.380 246.000 ;
        RECT 660.540 245.700 679.540 246.000 ;
        RECT 680.700 245.700 699.700 246.000 ;
        RECT 700.860 245.700 719.860 246.000 ;
        RECT 721.020 245.700 740.020 246.000 ;
        RECT 741.180 245.700 760.180 246.000 ;
        RECT 761.340 245.700 780.340 246.000 ;
        RECT 781.500 245.700 800.500 246.000 ;
        RECT 801.660 245.700 820.660 246.000 ;
        RECT 821.820 245.700 840.820 246.000 ;
        RECT 841.980 245.700 860.980 246.000 ;
        RECT 862.140 245.700 881.140 246.000 ;
        RECT 882.300 245.700 901.300 246.000 ;
        RECT 902.460 245.700 921.460 246.000 ;
        RECT 922.620 245.700 941.620 246.000 ;
        RECT 942.780 245.700 961.780 246.000 ;
        RECT 962.940 245.700 981.940 246.000 ;
        RECT 983.100 245.700 1002.100 246.000 ;
        RECT 1003.260 245.700 1022.260 246.000 ;
        RECT 1023.420 245.700 1042.420 246.000 ;
        RECT 1043.580 245.700 1062.580 246.000 ;
        RECT 1063.740 245.700 1082.740 246.000 ;
        RECT 1083.900 245.700 1087.940 246.000 ;
        RECT 14.700 4.300 1087.940 245.700 ;
        RECT 14.700 4.000 17.620 4.300 ;
        RECT 18.780 4.000 31.060 4.300 ;
        RECT 32.220 4.000 44.500 4.300 ;
        RECT 45.660 4.000 57.940 4.300 ;
        RECT 59.100 4.000 71.380 4.300 ;
        RECT 72.540 4.000 84.820 4.300 ;
        RECT 85.980 4.000 98.260 4.300 ;
        RECT 99.420 4.000 111.700 4.300 ;
        RECT 112.860 4.000 125.140 4.300 ;
        RECT 126.300 4.000 138.580 4.300 ;
        RECT 139.740 4.000 152.020 4.300 ;
        RECT 153.180 4.000 165.460 4.300 ;
        RECT 166.620 4.000 178.900 4.300 ;
        RECT 180.060 4.000 192.340 4.300 ;
        RECT 193.500 4.000 205.780 4.300 ;
        RECT 206.940 4.000 219.220 4.300 ;
        RECT 220.380 4.000 232.660 4.300 ;
        RECT 233.820 4.000 246.100 4.300 ;
        RECT 247.260 4.000 259.540 4.300 ;
        RECT 260.700 4.000 272.980 4.300 ;
        RECT 274.140 4.000 286.420 4.300 ;
        RECT 287.580 4.000 299.860 4.300 ;
        RECT 301.020 4.000 313.300 4.300 ;
        RECT 314.460 4.000 326.740 4.300 ;
        RECT 327.900 4.000 340.180 4.300 ;
        RECT 341.340 4.000 353.620 4.300 ;
        RECT 354.780 4.000 367.060 4.300 ;
        RECT 368.220 4.000 380.500 4.300 ;
        RECT 381.660 4.000 393.940 4.300 ;
        RECT 395.100 4.000 407.380 4.300 ;
        RECT 408.540 4.000 420.820 4.300 ;
        RECT 421.980 4.000 434.260 4.300 ;
        RECT 435.420 4.000 447.700 4.300 ;
        RECT 448.860 4.000 461.140 4.300 ;
        RECT 462.300 4.000 474.580 4.300 ;
        RECT 475.740 4.000 488.020 4.300 ;
        RECT 489.180 4.000 501.460 4.300 ;
        RECT 502.620 4.000 514.900 4.300 ;
        RECT 516.060 4.000 528.340 4.300 ;
        RECT 529.500 4.000 541.780 4.300 ;
        RECT 542.940 4.000 555.220 4.300 ;
        RECT 556.380 4.000 568.660 4.300 ;
        RECT 569.820 4.000 582.100 4.300 ;
        RECT 583.260 4.000 595.540 4.300 ;
        RECT 596.700 4.000 608.980 4.300 ;
        RECT 610.140 4.000 622.420 4.300 ;
        RECT 623.580 4.000 635.860 4.300 ;
        RECT 637.020 4.000 649.300 4.300 ;
        RECT 650.460 4.000 662.740 4.300 ;
        RECT 663.900 4.000 676.180 4.300 ;
        RECT 677.340 4.000 689.620 4.300 ;
        RECT 690.780 4.000 703.060 4.300 ;
        RECT 704.220 4.000 716.500 4.300 ;
        RECT 717.660 4.000 729.940 4.300 ;
        RECT 731.100 4.000 743.380 4.300 ;
        RECT 744.540 4.000 756.820 4.300 ;
        RECT 757.980 4.000 770.260 4.300 ;
        RECT 771.420 4.000 783.700 4.300 ;
        RECT 784.860 4.000 797.140 4.300 ;
        RECT 798.300 4.000 810.580 4.300 ;
        RECT 811.740 4.000 824.020 4.300 ;
        RECT 825.180 4.000 837.460 4.300 ;
        RECT 838.620 4.000 850.900 4.300 ;
        RECT 852.060 4.000 864.340 4.300 ;
        RECT 865.500 4.000 877.780 4.300 ;
        RECT 878.940 4.000 891.220 4.300 ;
        RECT 892.380 4.000 904.660 4.300 ;
        RECT 905.820 4.000 918.100 4.300 ;
        RECT 919.260 4.000 931.540 4.300 ;
        RECT 932.700 4.000 944.980 4.300 ;
        RECT 946.140 4.000 958.420 4.300 ;
        RECT 959.580 4.000 971.860 4.300 ;
        RECT 973.020 4.000 985.300 4.300 ;
        RECT 986.460 4.000 998.740 4.300 ;
        RECT 999.900 4.000 1012.180 4.300 ;
        RECT 1013.340 4.000 1025.620 4.300 ;
        RECT 1026.780 4.000 1039.060 4.300 ;
        RECT 1040.220 4.000 1052.500 4.300 ;
        RECT 1053.660 4.000 1065.940 4.300 ;
        RECT 1067.100 4.000 1079.380 4.300 ;
        RECT 1080.540 4.000 1087.940 4.300 ;
      LAYER Metal3 ;
        RECT 14.650 6.860 1087.990 231.420 ;
      LAYER Metal4 ;
        RECT 688.940 21.930 713.140 35.190 ;
        RECT 715.340 21.930 789.940 35.190 ;
        RECT 792.140 21.930 820.260 35.190 ;
  END
END ram_controller
END LIBRARY

