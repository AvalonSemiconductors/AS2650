magic
tech gf180mcuD
magscale 1 10
timestamp 1701086215
<< nwell >>
rect 1258 45824 218710 46342
rect 1258 44281 218710 45120
rect 1258 44256 132685 44281
rect 1258 43527 139448 43552
rect 1258 42688 218710 43527
rect 1258 41120 218710 41984
rect 1258 39552 218710 40416
rect 1258 37984 218710 38848
rect 1258 36416 218710 37280
rect 1258 34848 218710 35712
rect 1258 33280 218710 34144
rect 1258 31712 218710 32576
rect 1258 30983 107976 31008
rect 1258 30169 218710 30983
rect 1258 30144 95208 30169
rect 1258 29415 99800 29440
rect 1258 28576 218710 29415
rect 1258 27008 218710 27872
rect 1258 25440 218710 26304
rect 1258 23872 218710 24736
rect 1258 22304 218710 23168
rect 1258 20736 218710 21600
rect 1258 19168 218710 20032
rect 1258 17600 218710 18464
rect 1258 16032 218710 16896
rect 1258 14464 218710 15328
rect 1258 12896 218710 13760
rect 1258 11328 218710 12192
rect 1258 10599 156270 10624
rect 1258 9760 218710 10599
rect 1258 9031 135261 9056
rect 1258 8217 218710 9031
rect 1258 8192 132797 8217
rect 1258 7463 131453 7488
rect 1258 6649 218710 7463
rect 1258 6624 132797 6649
rect 1258 5895 136157 5920
rect 1258 5056 218710 5895
rect 1258 4327 151614 4352
rect 1258 3488 218710 4327
<< pwell >>
rect 1258 45120 218710 45824
rect 1258 43552 218710 44256
rect 1258 41984 218710 42688
rect 1258 40416 218710 41120
rect 1258 38848 218710 39552
rect 1258 37280 218710 37984
rect 1258 35712 218710 36416
rect 1258 34144 218710 34848
rect 1258 32576 218710 33280
rect 1258 31008 218710 31712
rect 1258 29440 218710 30144
rect 1258 27872 218710 28576
rect 1258 26304 218710 27008
rect 1258 24736 218710 25440
rect 1258 23168 218710 23872
rect 1258 21600 218710 22304
rect 1258 20032 218710 20736
rect 1258 18464 218710 19168
rect 1258 16896 218710 17600
rect 1258 15328 218710 16032
rect 1258 13760 218710 14464
rect 1258 12192 218710 12896
rect 1258 10624 218710 11328
rect 1258 9056 218710 9760
rect 1258 7488 218710 8192
rect 1258 5920 218710 6624
rect 1258 4352 218710 5056
rect 1258 3050 218710 3488
<< obsm1 >>
rect 1344 3076 218624 46450
<< metal2 >>
rect 2912 49200 3024 50000
rect 6944 49200 7056 50000
rect 10976 49200 11088 50000
rect 15008 49200 15120 50000
rect 19040 49200 19152 50000
rect 23072 49200 23184 50000
rect 27104 49200 27216 50000
rect 31136 49200 31248 50000
rect 35168 49200 35280 50000
rect 39200 49200 39312 50000
rect 43232 49200 43344 50000
rect 47264 49200 47376 50000
rect 51296 49200 51408 50000
rect 55328 49200 55440 50000
rect 59360 49200 59472 50000
rect 63392 49200 63504 50000
rect 67424 49200 67536 50000
rect 71456 49200 71568 50000
rect 75488 49200 75600 50000
rect 79520 49200 79632 50000
rect 83552 49200 83664 50000
rect 87584 49200 87696 50000
rect 91616 49200 91728 50000
rect 95648 49200 95760 50000
rect 99680 49200 99792 50000
rect 103712 49200 103824 50000
rect 107744 49200 107856 50000
rect 111776 49200 111888 50000
rect 115808 49200 115920 50000
rect 119840 49200 119952 50000
rect 123872 49200 123984 50000
rect 127904 49200 128016 50000
rect 131936 49200 132048 50000
rect 135968 49200 136080 50000
rect 140000 49200 140112 50000
rect 144032 49200 144144 50000
rect 148064 49200 148176 50000
rect 152096 49200 152208 50000
rect 156128 49200 156240 50000
rect 160160 49200 160272 50000
rect 164192 49200 164304 50000
rect 168224 49200 168336 50000
rect 172256 49200 172368 50000
rect 176288 49200 176400 50000
rect 180320 49200 180432 50000
rect 184352 49200 184464 50000
rect 188384 49200 188496 50000
rect 192416 49200 192528 50000
rect 196448 49200 196560 50000
rect 200480 49200 200592 50000
rect 204512 49200 204624 50000
rect 208544 49200 208656 50000
rect 212576 49200 212688 50000
rect 216608 49200 216720 50000
rect 3584 0 3696 800
rect 6272 0 6384 800
rect 8960 0 9072 800
rect 11648 0 11760 800
rect 14336 0 14448 800
rect 17024 0 17136 800
rect 19712 0 19824 800
rect 22400 0 22512 800
rect 25088 0 25200 800
rect 27776 0 27888 800
rect 30464 0 30576 800
rect 33152 0 33264 800
rect 35840 0 35952 800
rect 38528 0 38640 800
rect 41216 0 41328 800
rect 43904 0 44016 800
rect 46592 0 46704 800
rect 49280 0 49392 800
rect 51968 0 52080 800
rect 54656 0 54768 800
rect 57344 0 57456 800
rect 60032 0 60144 800
rect 62720 0 62832 800
rect 65408 0 65520 800
rect 68096 0 68208 800
rect 70784 0 70896 800
rect 73472 0 73584 800
rect 76160 0 76272 800
rect 78848 0 78960 800
rect 81536 0 81648 800
rect 84224 0 84336 800
rect 86912 0 87024 800
rect 89600 0 89712 800
rect 92288 0 92400 800
rect 94976 0 95088 800
rect 97664 0 97776 800
rect 100352 0 100464 800
rect 103040 0 103152 800
rect 105728 0 105840 800
rect 108416 0 108528 800
rect 111104 0 111216 800
rect 113792 0 113904 800
rect 116480 0 116592 800
rect 119168 0 119280 800
rect 121856 0 121968 800
rect 124544 0 124656 800
rect 127232 0 127344 800
rect 129920 0 130032 800
rect 132608 0 132720 800
rect 135296 0 135408 800
rect 137984 0 138096 800
rect 140672 0 140784 800
rect 143360 0 143472 800
rect 146048 0 146160 800
rect 148736 0 148848 800
rect 151424 0 151536 800
rect 154112 0 154224 800
rect 156800 0 156912 800
rect 159488 0 159600 800
rect 162176 0 162288 800
rect 164864 0 164976 800
rect 167552 0 167664 800
rect 170240 0 170352 800
rect 172928 0 173040 800
rect 175616 0 175728 800
rect 178304 0 178416 800
rect 180992 0 181104 800
rect 183680 0 183792 800
rect 186368 0 186480 800
rect 189056 0 189168 800
rect 191744 0 191856 800
rect 194432 0 194544 800
rect 197120 0 197232 800
rect 199808 0 199920 800
rect 202496 0 202608 800
rect 205184 0 205296 800
rect 207872 0 207984 800
rect 210560 0 210672 800
rect 213248 0 213360 800
rect 215936 0 216048 800
<< obsm2 >>
rect 3084 49140 6884 49200
rect 7116 49140 10916 49200
rect 11148 49140 14948 49200
rect 15180 49140 18980 49200
rect 19212 49140 23012 49200
rect 23244 49140 27044 49200
rect 27276 49140 31076 49200
rect 31308 49140 35108 49200
rect 35340 49140 39140 49200
rect 39372 49140 43172 49200
rect 43404 49140 47204 49200
rect 47436 49140 51236 49200
rect 51468 49140 55268 49200
rect 55500 49140 59300 49200
rect 59532 49140 63332 49200
rect 63564 49140 67364 49200
rect 67596 49140 71396 49200
rect 71628 49140 75428 49200
rect 75660 49140 79460 49200
rect 79692 49140 83492 49200
rect 83724 49140 87524 49200
rect 87756 49140 91556 49200
rect 91788 49140 95588 49200
rect 95820 49140 99620 49200
rect 99852 49140 103652 49200
rect 103884 49140 107684 49200
rect 107916 49140 111716 49200
rect 111948 49140 115748 49200
rect 115980 49140 119780 49200
rect 120012 49140 123812 49200
rect 124044 49140 127844 49200
rect 128076 49140 131876 49200
rect 132108 49140 135908 49200
rect 136140 49140 139940 49200
rect 140172 49140 143972 49200
rect 144204 49140 148004 49200
rect 148236 49140 152036 49200
rect 152268 49140 156068 49200
rect 156300 49140 160100 49200
rect 160332 49140 164132 49200
rect 164364 49140 168164 49200
rect 168396 49140 172196 49200
rect 172428 49140 176228 49200
rect 176460 49140 180260 49200
rect 180492 49140 184292 49200
rect 184524 49140 188324 49200
rect 188556 49140 192356 49200
rect 192588 49140 196388 49200
rect 196620 49140 200420 49200
rect 200652 49140 204452 49200
rect 204684 49140 208484 49200
rect 208716 49140 212516 49200
rect 212748 49140 216548 49200
rect 216780 49140 217588 49200
rect 2940 860 217588 49140
rect 2940 800 3524 860
rect 3756 800 6212 860
rect 6444 800 8900 860
rect 9132 800 11588 860
rect 11820 800 14276 860
rect 14508 800 16964 860
rect 17196 800 19652 860
rect 19884 800 22340 860
rect 22572 800 25028 860
rect 25260 800 27716 860
rect 27948 800 30404 860
rect 30636 800 33092 860
rect 33324 800 35780 860
rect 36012 800 38468 860
rect 38700 800 41156 860
rect 41388 800 43844 860
rect 44076 800 46532 860
rect 46764 800 49220 860
rect 49452 800 51908 860
rect 52140 800 54596 860
rect 54828 800 57284 860
rect 57516 800 59972 860
rect 60204 800 62660 860
rect 62892 800 65348 860
rect 65580 800 68036 860
rect 68268 800 70724 860
rect 70956 800 73412 860
rect 73644 800 76100 860
rect 76332 800 78788 860
rect 79020 800 81476 860
rect 81708 800 84164 860
rect 84396 800 86852 860
rect 87084 800 89540 860
rect 89772 800 92228 860
rect 92460 800 94916 860
rect 95148 800 97604 860
rect 97836 800 100292 860
rect 100524 800 102980 860
rect 103212 800 105668 860
rect 105900 800 108356 860
rect 108588 800 111044 860
rect 111276 800 113732 860
rect 113964 800 116420 860
rect 116652 800 119108 860
rect 119340 800 121796 860
rect 122028 800 124484 860
rect 124716 800 127172 860
rect 127404 800 129860 860
rect 130092 800 132548 860
rect 132780 800 135236 860
rect 135468 800 137924 860
rect 138156 800 140612 860
rect 140844 800 143300 860
rect 143532 800 145988 860
rect 146220 800 148676 860
rect 148908 800 151364 860
rect 151596 800 154052 860
rect 154284 800 156740 860
rect 156972 800 159428 860
rect 159660 800 162116 860
rect 162348 800 164804 860
rect 165036 800 167492 860
rect 167724 800 170180 860
rect 170412 800 172868 860
rect 173100 800 175556 860
rect 175788 800 178244 860
rect 178476 800 180932 860
rect 181164 800 183620 860
rect 183852 800 186308 860
rect 186540 800 188996 860
rect 189228 800 191684 860
rect 191916 800 194372 860
rect 194604 800 197060 860
rect 197292 800 199748 860
rect 199980 800 202436 860
rect 202668 800 205124 860
rect 205356 800 207812 860
rect 208044 800 210500 860
rect 210732 800 213188 860
rect 213420 800 215876 860
rect 216108 800 217588 860
<< obsm3 >>
rect 2930 1372 217598 46284
<< metal4 >>
rect 4448 3076 4768 46316
rect 19808 3076 20128 46316
rect 35168 3076 35488 46316
rect 50528 3076 50848 46316
rect 65888 3076 66208 46316
rect 81248 3076 81568 46316
rect 96608 3076 96928 46316
rect 111968 3076 112288 46316
rect 127328 3076 127648 46316
rect 142688 3076 143008 46316
rect 158048 3076 158368 46316
rect 173408 3076 173728 46316
rect 188768 3076 189088 46316
rect 204128 3076 204448 46316
<< obsm4 >>
rect 137788 4386 142628 7038
rect 143068 4386 157988 7038
rect 158428 4386 164052 7038
<< labels >>
rlabel metal2 s 27776 0 27888 800 6 A_all[0]
port 1 nsew signal output
rlabel metal2 s 30464 0 30576 800 6 A_all[1]
port 2 nsew signal output
rlabel metal2 s 33152 0 33264 800 6 A_all[2]
port 3 nsew signal output
rlabel metal2 s 35840 0 35952 800 6 A_all[3]
port 4 nsew signal output
rlabel metal2 s 38528 0 38640 800 6 A_all[4]
port 5 nsew signal output
rlabel metal2 s 41216 0 41328 800 6 A_all[5]
port 6 nsew signal output
rlabel metal2 s 43904 0 44016 800 6 A_all[6]
port 7 nsew signal output
rlabel metal2 s 46592 0 46704 800 6 A_all[7]
port 8 nsew signal output
rlabel metal2 s 49280 0 49392 800 6 A_all[8]
port 9 nsew signal output
rlabel metal2 s 3584 0 3696 800 6 CEN_all
port 10 nsew signal output
rlabel metal2 s 51968 0 52080 800 6 D_all[0]
port 11 nsew signal output
rlabel metal2 s 54656 0 54768 800 6 D_all[1]
port 12 nsew signal output
rlabel metal2 s 57344 0 57456 800 6 D_all[2]
port 13 nsew signal output
rlabel metal2 s 60032 0 60144 800 6 D_all[3]
port 14 nsew signal output
rlabel metal2 s 62720 0 62832 800 6 D_all[4]
port 15 nsew signal output
rlabel metal2 s 65408 0 65520 800 6 D_all[5]
port 16 nsew signal output
rlabel metal2 s 68096 0 68208 800 6 D_all[6]
port 17 nsew signal output
rlabel metal2 s 70784 0 70896 800 6 D_all[7]
port 18 nsew signal output
rlabel metal2 s 73472 0 73584 800 6 GWEN_0
port 19 nsew signal output
rlabel metal2 s 76160 0 76272 800 6 GWEN_1
port 20 nsew signal output
rlabel metal2 s 78848 0 78960 800 6 GWEN_2
port 21 nsew signal output
rlabel metal2 s 81536 0 81648 800 6 GWEN_3
port 22 nsew signal output
rlabel metal2 s 84224 0 84336 800 6 GWEN_4
port 23 nsew signal output
rlabel metal2 s 86912 0 87024 800 6 GWEN_5
port 24 nsew signal output
rlabel metal2 s 148064 49200 148176 50000 6 GWEN_6
port 25 nsew signal output
rlabel metal2 s 152096 49200 152208 50000 6 GWEN_7
port 26 nsew signal output
rlabel metal2 s 89600 0 89712 800 6 Q0[0]
port 27 nsew signal input
rlabel metal2 s 92288 0 92400 800 6 Q0[1]
port 28 nsew signal input
rlabel metal2 s 94976 0 95088 800 6 Q0[2]
port 29 nsew signal input
rlabel metal2 s 97664 0 97776 800 6 Q0[3]
port 30 nsew signal input
rlabel metal2 s 100352 0 100464 800 6 Q0[4]
port 31 nsew signal input
rlabel metal2 s 103040 0 103152 800 6 Q0[5]
port 32 nsew signal input
rlabel metal2 s 105728 0 105840 800 6 Q0[6]
port 33 nsew signal input
rlabel metal2 s 108416 0 108528 800 6 Q0[7]
port 34 nsew signal input
rlabel metal2 s 111104 0 111216 800 6 Q1[0]
port 35 nsew signal input
rlabel metal2 s 113792 0 113904 800 6 Q1[1]
port 36 nsew signal input
rlabel metal2 s 116480 0 116592 800 6 Q1[2]
port 37 nsew signal input
rlabel metal2 s 119168 0 119280 800 6 Q1[3]
port 38 nsew signal input
rlabel metal2 s 121856 0 121968 800 6 Q1[4]
port 39 nsew signal input
rlabel metal2 s 124544 0 124656 800 6 Q1[5]
port 40 nsew signal input
rlabel metal2 s 127232 0 127344 800 6 Q1[6]
port 41 nsew signal input
rlabel metal2 s 129920 0 130032 800 6 Q1[7]
port 42 nsew signal input
rlabel metal2 s 132608 0 132720 800 6 Q2[0]
port 43 nsew signal input
rlabel metal2 s 135296 0 135408 800 6 Q2[1]
port 44 nsew signal input
rlabel metal2 s 137984 0 138096 800 6 Q2[2]
port 45 nsew signal input
rlabel metal2 s 140672 0 140784 800 6 Q2[3]
port 46 nsew signal input
rlabel metal2 s 143360 0 143472 800 6 Q2[4]
port 47 nsew signal input
rlabel metal2 s 146048 0 146160 800 6 Q2[5]
port 48 nsew signal input
rlabel metal2 s 148736 0 148848 800 6 Q2[6]
port 49 nsew signal input
rlabel metal2 s 151424 0 151536 800 6 Q2[7]
port 50 nsew signal input
rlabel metal2 s 154112 0 154224 800 6 Q3[0]
port 51 nsew signal input
rlabel metal2 s 156800 0 156912 800 6 Q3[1]
port 52 nsew signal input
rlabel metal2 s 159488 0 159600 800 6 Q3[2]
port 53 nsew signal input
rlabel metal2 s 162176 0 162288 800 6 Q3[3]
port 54 nsew signal input
rlabel metal2 s 164864 0 164976 800 6 Q3[4]
port 55 nsew signal input
rlabel metal2 s 167552 0 167664 800 6 Q3[5]
port 56 nsew signal input
rlabel metal2 s 170240 0 170352 800 6 Q3[6]
port 57 nsew signal input
rlabel metal2 s 172928 0 173040 800 6 Q3[7]
port 58 nsew signal input
rlabel metal2 s 175616 0 175728 800 6 Q4[0]
port 59 nsew signal input
rlabel metal2 s 178304 0 178416 800 6 Q4[1]
port 60 nsew signal input
rlabel metal2 s 180992 0 181104 800 6 Q4[2]
port 61 nsew signal input
rlabel metal2 s 183680 0 183792 800 6 Q4[3]
port 62 nsew signal input
rlabel metal2 s 186368 0 186480 800 6 Q4[4]
port 63 nsew signal input
rlabel metal2 s 189056 0 189168 800 6 Q4[5]
port 64 nsew signal input
rlabel metal2 s 191744 0 191856 800 6 Q4[6]
port 65 nsew signal input
rlabel metal2 s 194432 0 194544 800 6 Q4[7]
port 66 nsew signal input
rlabel metal2 s 197120 0 197232 800 6 Q5[0]
port 67 nsew signal input
rlabel metal2 s 199808 0 199920 800 6 Q5[1]
port 68 nsew signal input
rlabel metal2 s 202496 0 202608 800 6 Q5[2]
port 69 nsew signal input
rlabel metal2 s 205184 0 205296 800 6 Q5[3]
port 70 nsew signal input
rlabel metal2 s 207872 0 207984 800 6 Q5[4]
port 71 nsew signal input
rlabel metal2 s 210560 0 210672 800 6 Q5[5]
port 72 nsew signal input
rlabel metal2 s 213248 0 213360 800 6 Q5[6]
port 73 nsew signal input
rlabel metal2 s 215936 0 216048 800 6 Q5[7]
port 74 nsew signal input
rlabel metal2 s 156128 49200 156240 50000 6 Q6[0]
port 75 nsew signal input
rlabel metal2 s 160160 49200 160272 50000 6 Q6[1]
port 76 nsew signal input
rlabel metal2 s 164192 49200 164304 50000 6 Q6[2]
port 77 nsew signal input
rlabel metal2 s 168224 49200 168336 50000 6 Q6[3]
port 78 nsew signal input
rlabel metal2 s 172256 49200 172368 50000 6 Q6[4]
port 79 nsew signal input
rlabel metal2 s 176288 49200 176400 50000 6 Q6[5]
port 80 nsew signal input
rlabel metal2 s 180320 49200 180432 50000 6 Q6[6]
port 81 nsew signal input
rlabel metal2 s 184352 49200 184464 50000 6 Q6[7]
port 82 nsew signal input
rlabel metal2 s 188384 49200 188496 50000 6 Q7[0]
port 83 nsew signal input
rlabel metal2 s 192416 49200 192528 50000 6 Q7[1]
port 84 nsew signal input
rlabel metal2 s 196448 49200 196560 50000 6 Q7[2]
port 85 nsew signal input
rlabel metal2 s 200480 49200 200592 50000 6 Q7[3]
port 86 nsew signal input
rlabel metal2 s 204512 49200 204624 50000 6 Q7[4]
port 87 nsew signal input
rlabel metal2 s 208544 49200 208656 50000 6 Q7[5]
port 88 nsew signal input
rlabel metal2 s 212576 49200 212688 50000 6 Q7[6]
port 89 nsew signal input
rlabel metal2 s 216608 49200 216720 50000 6 Q7[7]
port 90 nsew signal input
rlabel metal2 s 6272 0 6384 800 6 WEN_all[0]
port 91 nsew signal output
rlabel metal2 s 8960 0 9072 800 6 WEN_all[1]
port 92 nsew signal output
rlabel metal2 s 11648 0 11760 800 6 WEN_all[2]
port 93 nsew signal output
rlabel metal2 s 14336 0 14448 800 6 WEN_all[3]
port 94 nsew signal output
rlabel metal2 s 17024 0 17136 800 6 WEN_all[4]
port 95 nsew signal output
rlabel metal2 s 19712 0 19824 800 6 WEN_all[5]
port 96 nsew signal output
rlabel metal2 s 22400 0 22512 800 6 WEN_all[6]
port 97 nsew signal output
rlabel metal2 s 25088 0 25200 800 6 WEN_all[7]
port 98 nsew signal output
rlabel metal2 s 10976 49200 11088 50000 6 WEb_ram
port 99 nsew signal input
rlabel metal2 s 15008 49200 15120 50000 6 bus_in[0]
port 100 nsew signal input
rlabel metal2 s 19040 49200 19152 50000 6 bus_in[1]
port 101 nsew signal input
rlabel metal2 s 23072 49200 23184 50000 6 bus_in[2]
port 102 nsew signal input
rlabel metal2 s 27104 49200 27216 50000 6 bus_in[3]
port 103 nsew signal input
rlabel metal2 s 31136 49200 31248 50000 6 bus_in[4]
port 104 nsew signal input
rlabel metal2 s 35168 49200 35280 50000 6 bus_in[5]
port 105 nsew signal input
rlabel metal2 s 39200 49200 39312 50000 6 bus_in[6]
port 106 nsew signal input
rlabel metal2 s 43232 49200 43344 50000 6 bus_in[7]
port 107 nsew signal input
rlabel metal2 s 47264 49200 47376 50000 6 bus_out[0]
port 108 nsew signal output
rlabel metal2 s 51296 49200 51408 50000 6 bus_out[1]
port 109 nsew signal output
rlabel metal2 s 55328 49200 55440 50000 6 bus_out[2]
port 110 nsew signal output
rlabel metal2 s 59360 49200 59472 50000 6 bus_out[3]
port 111 nsew signal output
rlabel metal2 s 63392 49200 63504 50000 6 bus_out[4]
port 112 nsew signal output
rlabel metal2 s 67424 49200 67536 50000 6 bus_out[5]
port 113 nsew signal output
rlabel metal2 s 71456 49200 71568 50000 6 bus_out[6]
port 114 nsew signal output
rlabel metal2 s 75488 49200 75600 50000 6 bus_out[7]
port 115 nsew signal output
rlabel metal2 s 79520 49200 79632 50000 6 ram_enabled
port 116 nsew signal input
rlabel metal2 s 83552 49200 83664 50000 6 requested_addr[0]
port 117 nsew signal input
rlabel metal2 s 123872 49200 123984 50000 6 requested_addr[10]
port 118 nsew signal input
rlabel metal2 s 127904 49200 128016 50000 6 requested_addr[11]
port 119 nsew signal input
rlabel metal2 s 131936 49200 132048 50000 6 requested_addr[12]
port 120 nsew signal input
rlabel metal2 s 135968 49200 136080 50000 6 requested_addr[13]
port 121 nsew signal input
rlabel metal2 s 140000 49200 140112 50000 6 requested_addr[14]
port 122 nsew signal input
rlabel metal2 s 144032 49200 144144 50000 6 requested_addr[15]
port 123 nsew signal input
rlabel metal2 s 87584 49200 87696 50000 6 requested_addr[1]
port 124 nsew signal input
rlabel metal2 s 91616 49200 91728 50000 6 requested_addr[2]
port 125 nsew signal input
rlabel metal2 s 95648 49200 95760 50000 6 requested_addr[3]
port 126 nsew signal input
rlabel metal2 s 99680 49200 99792 50000 6 requested_addr[4]
port 127 nsew signal input
rlabel metal2 s 103712 49200 103824 50000 6 requested_addr[5]
port 128 nsew signal input
rlabel metal2 s 107744 49200 107856 50000 6 requested_addr[6]
port 129 nsew signal input
rlabel metal2 s 111776 49200 111888 50000 6 requested_addr[7]
port 130 nsew signal input
rlabel metal2 s 115808 49200 115920 50000 6 requested_addr[8]
port 131 nsew signal input
rlabel metal2 s 119840 49200 119952 50000 6 requested_addr[9]
port 132 nsew signal input
rlabel metal2 s 6944 49200 7056 50000 6 rst
port 133 nsew signal input
rlabel metal4 s 4448 3076 4768 46316 6 vdd
port 134 nsew power bidirectional
rlabel metal4 s 35168 3076 35488 46316 6 vdd
port 134 nsew power bidirectional
rlabel metal4 s 65888 3076 66208 46316 6 vdd
port 134 nsew power bidirectional
rlabel metal4 s 96608 3076 96928 46316 6 vdd
port 134 nsew power bidirectional
rlabel metal4 s 127328 3076 127648 46316 6 vdd
port 134 nsew power bidirectional
rlabel metal4 s 158048 3076 158368 46316 6 vdd
port 134 nsew power bidirectional
rlabel metal4 s 188768 3076 189088 46316 6 vdd
port 134 nsew power bidirectional
rlabel metal4 s 19808 3076 20128 46316 6 vss
port 135 nsew ground bidirectional
rlabel metal4 s 50528 3076 50848 46316 6 vss
port 135 nsew ground bidirectional
rlabel metal4 s 81248 3076 81568 46316 6 vss
port 135 nsew ground bidirectional
rlabel metal4 s 111968 3076 112288 46316 6 vss
port 135 nsew ground bidirectional
rlabel metal4 s 142688 3076 143008 46316 6 vss
port 135 nsew ground bidirectional
rlabel metal4 s 173408 3076 173728 46316 6 vss
port 135 nsew ground bidirectional
rlabel metal4 s 204128 3076 204448 46316 6 vss
port 135 nsew ground bidirectional
rlabel metal2 s 2912 49200 3024 50000 6 wb_clk_i
port 136 nsew signal input
<< properties >>
string FIXED_BBOX 0 0 220000 50000
string LEFclass BLOCK
string LEFview TRUE
string GDS_END 1398572
string GDS_FILE /run/media/tholin/fbc90f8f-67e9-406d-9872-54f02ad6a2d8/AS2650/openlane/ram_controller/runs/23_11_27_12_52/results/signoff/ram_controller.magic.gds
string GDS_START 175762
<< end >>

