magic
tech gf180mcuD
magscale 1 10
timestamp 1700515028
<< metal1 >>
rect 38770 56590 38782 56642
rect 38834 56639 38846 56642
rect 39330 56639 39342 56642
rect 38834 56593 39342 56639
rect 38834 56590 38846 56593
rect 39330 56590 39342 56593
rect 39394 56639 39406 56642
rect 40114 56639 40126 56642
rect 39394 56593 40126 56639
rect 39394 56590 39406 56593
rect 40114 56590 40126 56593
rect 40178 56590 40190 56642
rect 1344 56474 58576 56508
rect 1344 56422 19838 56474
rect 19890 56422 19942 56474
rect 19994 56422 20046 56474
rect 20098 56422 50558 56474
rect 50610 56422 50662 56474
rect 50714 56422 50766 56474
rect 50818 56422 58576 56474
rect 1344 56388 58576 56422
rect 5070 56306 5122 56318
rect 5070 56242 5122 56254
rect 7422 56306 7474 56318
rect 7422 56242 7474 56254
rect 7646 56306 7698 56318
rect 7646 56242 7698 56254
rect 9662 56306 9714 56318
rect 9662 56242 9714 56254
rect 9886 56306 9938 56318
rect 9886 56242 9938 56254
rect 11902 56306 11954 56318
rect 11902 56242 11954 56254
rect 12126 56306 12178 56318
rect 12126 56242 12178 56254
rect 14142 56306 14194 56318
rect 14142 56242 14194 56254
rect 16494 56306 16546 56318
rect 16494 56242 16546 56254
rect 16942 56306 16994 56318
rect 16942 56242 16994 56254
rect 18622 56306 18674 56318
rect 18622 56242 18674 56254
rect 18846 56306 18898 56318
rect 18846 56242 18898 56254
rect 20302 56306 20354 56318
rect 20302 56242 20354 56254
rect 23102 56306 23154 56318
rect 23102 56242 23154 56254
rect 25342 56306 25394 56318
rect 25342 56242 25394 56254
rect 27918 56306 27970 56318
rect 27918 56242 27970 56254
rect 29822 56306 29874 56318
rect 29822 56242 29874 56254
rect 31726 56306 31778 56318
rect 31726 56242 31778 56254
rect 34302 56306 34354 56318
rect 34302 56242 34354 56254
rect 36542 56306 36594 56318
rect 36542 56242 36594 56254
rect 39342 56306 39394 56318
rect 39342 56242 39394 56254
rect 41470 56306 41522 56318
rect 41470 56242 41522 56254
rect 44606 56306 44658 56318
rect 44606 56242 44658 56254
rect 48974 56306 49026 56318
rect 48974 56242 49026 56254
rect 52222 56306 52274 56318
rect 52222 56242 52274 56254
rect 56030 56306 56082 56318
rect 56030 56242 56082 56254
rect 2046 56194 2098 56206
rect 2046 56130 2098 56142
rect 2382 56194 2434 56206
rect 2382 56130 2434 56142
rect 5518 56194 5570 56206
rect 5518 56130 5570 56142
rect 5854 56194 5906 56206
rect 14366 56194 14418 56206
rect 21086 56194 21138 56206
rect 7970 56142 7982 56194
rect 8034 56142 8046 56194
rect 10210 56142 10222 56194
rect 10274 56142 10286 56194
rect 12450 56142 12462 56194
rect 12514 56142 12526 56194
rect 17266 56142 17278 56194
rect 17330 56142 17342 56194
rect 19170 56142 19182 56194
rect 19234 56142 19246 56194
rect 5854 56130 5906 56142
rect 14366 56130 14418 56142
rect 21086 56130 21138 56142
rect 21422 56194 21474 56206
rect 21422 56130 21474 56142
rect 23326 56194 23378 56206
rect 23326 56130 23378 56142
rect 25566 56194 25618 56206
rect 25566 56130 25618 56142
rect 28366 56194 28418 56206
rect 28366 56130 28418 56142
rect 30046 56194 30098 56206
rect 30046 56130 30098 56142
rect 32286 56194 32338 56206
rect 32286 56130 32338 56142
rect 32622 56194 32674 56206
rect 32622 56130 32674 56142
rect 34526 56194 34578 56206
rect 34526 56130 34578 56142
rect 34862 56194 34914 56206
rect 34862 56130 34914 56142
rect 36766 56194 36818 56206
rect 36766 56130 36818 56142
rect 37102 56194 37154 56206
rect 37102 56130 37154 56142
rect 39790 56194 39842 56206
rect 39790 56130 39842 56142
rect 40126 56194 40178 56206
rect 40126 56130 40178 56142
rect 1710 56082 1762 56094
rect 47742 56082 47794 56094
rect 54574 56082 54626 56094
rect 2594 56030 2606 56082
rect 2658 56030 2670 56082
rect 14578 56030 14590 56082
rect 14642 56030 14654 56082
rect 23538 56030 23550 56082
rect 23602 56030 23614 56082
rect 25778 56030 25790 56082
rect 25842 56030 25854 56082
rect 28578 56030 28590 56082
rect 28642 56030 28654 56082
rect 30258 56030 30270 56082
rect 30322 56030 30334 56082
rect 40450 56030 40462 56082
rect 40514 56030 40526 56082
rect 43698 56030 43710 56082
rect 43762 56030 43774 56082
rect 47954 56030 47966 56082
rect 48018 56030 48030 56082
rect 51202 56030 51214 56082
rect 51266 56030 51278 56082
rect 55010 56030 55022 56082
rect 55074 56030 55086 56082
rect 1710 56018 1762 56030
rect 47742 56018 47794 56030
rect 54574 56018 54626 56030
rect 3166 55970 3218 55982
rect 3166 55906 3218 55918
rect 37998 55970 38050 55982
rect 37998 55906 38050 55918
rect 38894 55970 38946 55982
rect 38894 55906 38946 55918
rect 1344 55690 58576 55724
rect 1344 55638 4478 55690
rect 4530 55638 4582 55690
rect 4634 55638 4686 55690
rect 4738 55638 35198 55690
rect 35250 55638 35302 55690
rect 35354 55638 35406 55690
rect 35458 55638 58576 55690
rect 1344 55604 58576 55638
rect 2158 55410 2210 55422
rect 39230 55410 39282 55422
rect 46734 55410 46786 55422
rect 16370 55358 16382 55410
rect 16434 55358 16446 55410
rect 20514 55358 20526 55410
rect 20578 55358 20590 55410
rect 32050 55358 32062 55410
rect 32114 55358 32126 55410
rect 36418 55358 36430 55410
rect 36482 55358 36494 55410
rect 43138 55358 43150 55410
rect 43202 55358 43214 55410
rect 2158 55346 2210 55358
rect 39230 55346 39282 55358
rect 46734 55346 46786 55358
rect 53678 55410 53730 55422
rect 56690 55358 56702 55410
rect 56754 55358 56766 55410
rect 53678 55346 53730 55358
rect 16830 55298 16882 55310
rect 21422 55298 21474 55310
rect 13570 55246 13582 55298
rect 13634 55246 13646 55298
rect 17714 55246 17726 55298
rect 17778 55246 17790 55298
rect 16830 55234 16882 55246
rect 21422 55234 21474 55246
rect 22990 55298 23042 55310
rect 22990 55234 23042 55246
rect 25342 55298 25394 55310
rect 25342 55234 25394 55246
rect 27694 55298 27746 55310
rect 33182 55298 33234 55310
rect 29250 55246 29262 55298
rect 29314 55246 29326 55298
rect 32610 55246 32622 55298
rect 32674 55246 32686 55298
rect 33618 55246 33630 55298
rect 33682 55246 33694 55298
rect 37090 55246 37102 55298
rect 37154 55246 37166 55298
rect 40338 55246 40350 55298
rect 40402 55246 40414 55298
rect 45714 55246 45726 55298
rect 45778 55246 45790 55298
rect 52658 55246 52670 55298
rect 52722 55246 52734 55298
rect 55570 55246 55582 55298
rect 55634 55246 55646 55298
rect 27694 55234 27746 55246
rect 33182 55234 33234 55246
rect 11790 55186 11842 55198
rect 14242 55134 14254 55186
rect 14306 55134 14318 55186
rect 18386 55134 18398 55186
rect 18450 55134 18462 55186
rect 29922 55134 29934 55186
rect 29986 55134 29998 55186
rect 34290 55134 34302 55186
rect 34354 55134 34366 55186
rect 37314 55134 37326 55186
rect 37378 55134 37390 55186
rect 41010 55134 41022 55186
rect 41074 55134 41086 55186
rect 11790 55122 11842 55134
rect 11902 55074 11954 55086
rect 11902 55010 11954 55022
rect 22878 55074 22930 55086
rect 22878 55010 22930 55022
rect 25230 55074 25282 55086
rect 25230 55010 25282 55022
rect 27582 55074 27634 55086
rect 27582 55010 27634 55022
rect 32622 55074 32674 55086
rect 32622 55010 32674 55022
rect 37774 55074 37826 55086
rect 38558 55074 38610 55086
rect 38210 55022 38222 55074
rect 38274 55022 38286 55074
rect 37774 55010 37826 55022
rect 38558 55010 38610 55022
rect 39118 55074 39170 55086
rect 39118 55010 39170 55022
rect 39902 55074 39954 55086
rect 39902 55010 39954 55022
rect 43598 55074 43650 55086
rect 43598 55010 43650 55022
rect 45390 55074 45442 55086
rect 45390 55010 45442 55022
rect 50878 55074 50930 55086
rect 50878 55010 50930 55022
rect 52110 55074 52162 55086
rect 52110 55010 52162 55022
rect 1344 54906 58576 54940
rect 1344 54854 19838 54906
rect 19890 54854 19942 54906
rect 19994 54854 20046 54906
rect 20098 54854 50558 54906
rect 50610 54854 50662 54906
rect 50714 54854 50766 54906
rect 50818 54854 58576 54906
rect 1344 54820 58576 54854
rect 12462 54738 12514 54750
rect 12462 54674 12514 54686
rect 14814 54738 14866 54750
rect 14814 54674 14866 54686
rect 15822 54738 15874 54750
rect 15822 54674 15874 54686
rect 17614 54738 17666 54750
rect 17614 54674 17666 54686
rect 18510 54738 18562 54750
rect 18510 54674 18562 54686
rect 29934 54738 29986 54750
rect 29934 54674 29986 54686
rect 33966 54738 34018 54750
rect 33966 54674 34018 54686
rect 36430 54738 36482 54750
rect 36430 54674 36482 54686
rect 40350 54738 40402 54750
rect 40350 54674 40402 54686
rect 40910 54738 40962 54750
rect 40910 54674 40962 54686
rect 2046 54626 2098 54638
rect 15262 54626 15314 54638
rect 12786 54574 12798 54626
rect 12850 54574 12862 54626
rect 13234 54574 13246 54626
rect 13298 54574 13310 54626
rect 2046 54562 2098 54574
rect 15262 54562 15314 54574
rect 18734 54626 18786 54638
rect 18734 54562 18786 54574
rect 29150 54626 29202 54638
rect 29150 54562 29202 54574
rect 29486 54626 29538 54638
rect 29486 54562 29538 54574
rect 31838 54626 31890 54638
rect 31838 54562 31890 54574
rect 34750 54626 34802 54638
rect 34750 54562 34802 54574
rect 36654 54626 36706 54638
rect 41694 54626 41746 54638
rect 38882 54574 38894 54626
rect 38946 54574 38958 54626
rect 36654 54562 36706 54574
rect 41694 54562 41746 54574
rect 1710 54514 1762 54526
rect 14590 54514 14642 54526
rect 13682 54462 13694 54514
rect 13746 54462 13758 54514
rect 1710 54450 1762 54462
rect 14590 54450 14642 54462
rect 15038 54514 15090 54526
rect 15038 54450 15090 54462
rect 15710 54514 15762 54526
rect 15710 54450 15762 54462
rect 15934 54514 15986 54526
rect 15934 54450 15986 54462
rect 16382 54514 16434 54526
rect 16382 54450 16434 54462
rect 17278 54514 17330 54526
rect 17278 54450 17330 54462
rect 17726 54514 17778 54526
rect 17726 54450 17778 54462
rect 17838 54514 17890 54526
rect 17838 54450 17890 54462
rect 18286 54514 18338 54526
rect 18286 54450 18338 54462
rect 18398 54514 18450 54526
rect 28814 54514 28866 54526
rect 21074 54462 21086 54514
rect 21138 54462 21150 54514
rect 25330 54462 25342 54514
rect 25394 54462 25406 54514
rect 18398 54450 18450 54462
rect 28814 54450 28866 54462
rect 29822 54514 29874 54526
rect 33182 54514 33234 54526
rect 38558 54514 38610 54526
rect 41358 54514 41410 54526
rect 30034 54462 30046 54514
rect 30098 54462 30110 54514
rect 30594 54462 30606 54514
rect 30658 54462 30670 54514
rect 33394 54462 33406 54514
rect 33458 54462 33470 54514
rect 33954 54462 33966 54514
rect 34018 54462 34030 54514
rect 41010 54462 41022 54514
rect 41074 54462 41086 54514
rect 29822 54450 29874 54462
rect 33182 54450 33234 54462
rect 38558 54450 38610 54462
rect 41358 54450 41410 54462
rect 2494 54402 2546 54414
rect 32510 54402 32562 54414
rect 38222 54402 38274 54414
rect 13794 54350 13806 54402
rect 13858 54350 13870 54402
rect 21746 54350 21758 54402
rect 21810 54350 21822 54402
rect 23874 54350 23886 54402
rect 23938 54350 23950 54402
rect 26002 54350 26014 54402
rect 26066 54350 26078 54402
rect 28130 54350 28142 54402
rect 28194 54350 28206 54402
rect 31714 54350 31726 54402
rect 31778 54350 31790 54402
rect 34402 54350 34414 54402
rect 34466 54350 34478 54402
rect 36306 54350 36318 54402
rect 36370 54350 36382 54402
rect 2494 54338 2546 54350
rect 32510 54338 32562 54350
rect 38222 54338 38274 54350
rect 55246 54402 55298 54414
rect 55246 54338 55298 54350
rect 32062 54290 32114 54302
rect 30370 54238 30382 54290
rect 30434 54238 30446 54290
rect 32062 54226 32114 54238
rect 33630 54290 33682 54302
rect 33630 54226 33682 54238
rect 41246 54290 41298 54302
rect 41246 54226 41298 54238
rect 1344 54122 58576 54156
rect 1344 54070 4478 54122
rect 4530 54070 4582 54122
rect 4634 54070 4686 54122
rect 4738 54070 35198 54122
rect 35250 54070 35302 54122
rect 35354 54070 35406 54122
rect 35458 54070 58576 54122
rect 1344 54036 58576 54070
rect 40910 53954 40962 53966
rect 40910 53890 40962 53902
rect 23662 53842 23714 53854
rect 23662 53778 23714 53790
rect 29262 53842 29314 53854
rect 29262 53778 29314 53790
rect 41022 53842 41074 53854
rect 42130 53790 42142 53842
rect 42194 53790 42206 53842
rect 41022 53778 41074 53790
rect 22430 53730 22482 53742
rect 22430 53666 22482 53678
rect 22654 53730 22706 53742
rect 22654 53666 22706 53678
rect 22878 53730 22930 53742
rect 22878 53666 22930 53678
rect 23774 53730 23826 53742
rect 23774 53666 23826 53678
rect 24558 53730 24610 53742
rect 33058 53678 33070 53730
rect 33122 53678 33134 53730
rect 38322 53678 38334 53730
rect 38386 53678 38398 53730
rect 41234 53678 41246 53730
rect 41298 53678 41310 53730
rect 24558 53666 24610 53678
rect 22318 53618 22370 53630
rect 22318 53554 22370 53566
rect 25006 53618 25058 53630
rect 25006 53554 25058 53566
rect 25230 53618 25282 53630
rect 25230 53554 25282 53566
rect 26350 53618 26402 53630
rect 26350 53554 26402 53566
rect 32622 53618 32674 53630
rect 32622 53554 32674 53566
rect 33294 53618 33346 53630
rect 33294 53554 33346 53566
rect 37774 53618 37826 53630
rect 37774 53554 37826 53566
rect 38782 53618 38834 53630
rect 38782 53554 38834 53566
rect 39118 53618 39170 53630
rect 39118 53554 39170 53566
rect 42478 53618 42530 53630
rect 42478 53554 42530 53566
rect 10446 53506 10498 53518
rect 10446 53442 10498 53454
rect 11566 53506 11618 53518
rect 11566 53442 11618 53454
rect 15486 53506 15538 53518
rect 15486 53442 15538 53454
rect 16046 53506 16098 53518
rect 16046 53442 16098 53454
rect 16382 53506 16434 53518
rect 18174 53506 18226 53518
rect 16706 53454 16718 53506
rect 16770 53454 16782 53506
rect 16382 53442 16434 53454
rect 18174 53442 18226 53454
rect 21982 53506 22034 53518
rect 21982 53442 22034 53454
rect 23550 53506 23602 53518
rect 23550 53442 23602 53454
rect 23998 53506 24050 53518
rect 23998 53442 24050 53454
rect 24894 53506 24946 53518
rect 24894 53442 24946 53454
rect 25678 53506 25730 53518
rect 25678 53442 25730 53454
rect 26238 53506 26290 53518
rect 26238 53442 26290 53454
rect 26462 53506 26514 53518
rect 26462 53442 26514 53454
rect 26686 53506 26738 53518
rect 42254 53506 42306 53518
rect 38098 53454 38110 53506
rect 38162 53454 38174 53506
rect 26686 53442 26738 53454
rect 42254 53442 42306 53454
rect 1344 53338 58576 53372
rect 1344 53286 19838 53338
rect 19890 53286 19942 53338
rect 19994 53286 20046 53338
rect 20098 53286 50558 53338
rect 50610 53286 50662 53338
rect 50714 53286 50766 53338
rect 50818 53286 58576 53338
rect 1344 53252 58576 53286
rect 12798 53170 12850 53182
rect 12798 53106 12850 53118
rect 23438 53170 23490 53182
rect 23438 53106 23490 53118
rect 29262 53170 29314 53182
rect 29262 53106 29314 53118
rect 32062 53170 32114 53182
rect 32062 53106 32114 53118
rect 33966 53170 34018 53182
rect 33966 53106 34018 53118
rect 38446 53170 38498 53182
rect 38446 53106 38498 53118
rect 41022 53170 41074 53182
rect 41022 53106 41074 53118
rect 2046 53058 2098 53070
rect 2046 52994 2098 53006
rect 9886 53058 9938 53070
rect 9886 52994 9938 53006
rect 10558 53058 10610 53070
rect 10558 52994 10610 53006
rect 12014 53058 12066 53070
rect 12014 52994 12066 53006
rect 12350 53058 12402 53070
rect 12350 52994 12402 53006
rect 22766 53058 22818 53070
rect 29710 53058 29762 53070
rect 26674 53006 26686 53058
rect 26738 53006 26750 53058
rect 22766 52994 22818 53006
rect 29710 52994 29762 53006
rect 30046 53058 30098 53070
rect 32286 53058 32338 53070
rect 30258 53006 30270 53058
rect 30322 53006 30334 53058
rect 30046 52994 30098 53006
rect 32286 52994 32338 53006
rect 36654 53058 36706 53070
rect 36654 52994 36706 53006
rect 36766 53058 36818 53070
rect 36766 52994 36818 53006
rect 1710 52946 1762 52958
rect 10222 52946 10274 52958
rect 7970 52894 7982 52946
rect 8034 52894 8046 52946
rect 8754 52894 8766 52946
rect 8818 52894 8830 52946
rect 1710 52882 1762 52894
rect 10222 52882 10274 52894
rect 10670 52946 10722 52958
rect 10670 52882 10722 52894
rect 10894 52946 10946 52958
rect 18062 52946 18114 52958
rect 11330 52894 11342 52946
rect 11394 52894 11406 52946
rect 10894 52882 10946 52894
rect 18062 52882 18114 52894
rect 18398 52946 18450 52958
rect 18398 52882 18450 52894
rect 18510 52946 18562 52958
rect 18510 52882 18562 52894
rect 22430 52946 22482 52958
rect 22430 52882 22482 52894
rect 22990 52946 23042 52958
rect 22990 52882 23042 52894
rect 25454 52946 25506 52958
rect 25454 52882 25506 52894
rect 25902 52946 25954 52958
rect 25902 52882 25954 52894
rect 26126 52946 26178 52958
rect 26126 52882 26178 52894
rect 27022 52946 27074 52958
rect 27022 52882 27074 52894
rect 30494 52946 30546 52958
rect 33182 52946 33234 52958
rect 33630 52946 33682 52958
rect 36542 52946 36594 52958
rect 37774 52946 37826 52958
rect 30818 52894 30830 52946
rect 30882 52894 30894 52946
rect 33394 52894 33406 52946
rect 33458 52894 33470 52946
rect 33954 52894 33966 52946
rect 34018 52894 34030 52946
rect 36978 52894 36990 52946
rect 37042 52894 37054 52946
rect 37986 52894 37998 52946
rect 38050 52894 38062 52946
rect 41906 52894 41918 52946
rect 41970 52894 41982 52946
rect 42690 52894 42702 52946
rect 42754 52894 42766 52946
rect 30494 52882 30546 52894
rect 33182 52882 33234 52894
rect 33630 52882 33682 52894
rect 36542 52882 36594 52894
rect 37774 52882 37826 52894
rect 2494 52834 2546 52846
rect 15374 52834 15426 52846
rect 5842 52782 5854 52834
rect 5906 52782 5918 52834
rect 2494 52770 2546 52782
rect 15374 52770 15426 52782
rect 18174 52834 18226 52846
rect 18174 52770 18226 52782
rect 19070 52834 19122 52846
rect 19070 52770 19122 52782
rect 22542 52834 22594 52846
rect 22542 52770 22594 52782
rect 26014 52834 26066 52846
rect 26014 52770 26066 52782
rect 27470 52834 27522 52846
rect 27470 52770 27522 52782
rect 30158 52834 30210 52846
rect 37662 52834 37714 52846
rect 31938 52782 31950 52834
rect 32002 52782 32014 52834
rect 30158 52770 30210 52782
rect 37662 52770 37714 52782
rect 41582 52834 41634 52846
rect 44818 52782 44830 52834
rect 44882 52782 44894 52834
rect 41582 52770 41634 52782
rect 11006 52722 11058 52734
rect 11006 52658 11058 52670
rect 29598 52722 29650 52734
rect 29598 52658 29650 52670
rect 37438 52722 37490 52734
rect 41010 52670 41022 52722
rect 41074 52719 41086 52722
rect 41458 52719 41470 52722
rect 41074 52673 41470 52719
rect 41074 52670 41086 52673
rect 41458 52670 41470 52673
rect 41522 52670 41534 52722
rect 37438 52658 37490 52670
rect 1344 52554 58576 52588
rect 1344 52502 4478 52554
rect 4530 52502 4582 52554
rect 4634 52502 4686 52554
rect 4738 52502 35198 52554
rect 35250 52502 35302 52554
rect 35354 52502 35406 52554
rect 35458 52502 58576 52554
rect 1344 52468 58576 52502
rect 10446 52386 10498 52398
rect 41694 52386 41746 52398
rect 11666 52334 11678 52386
rect 11730 52334 11742 52386
rect 12002 52334 12014 52386
rect 12066 52383 12078 52386
rect 13010 52383 13022 52386
rect 12066 52337 13022 52383
rect 12066 52334 12078 52337
rect 13010 52334 13022 52337
rect 13074 52334 13086 52386
rect 10446 52322 10498 52334
rect 41694 52322 41746 52334
rect 12798 52274 12850 52286
rect 32846 52274 32898 52286
rect 17826 52222 17838 52274
rect 17890 52222 17902 52274
rect 19954 52222 19966 52274
rect 20018 52222 20030 52274
rect 30146 52222 30158 52274
rect 30210 52222 30222 52274
rect 32274 52222 32286 52274
rect 32338 52222 32350 52274
rect 34178 52222 34190 52274
rect 34242 52222 34254 52274
rect 36306 52222 36318 52274
rect 36370 52222 36382 52274
rect 38658 52222 38670 52274
rect 38722 52222 38734 52274
rect 42690 52222 42702 52274
rect 42754 52222 42766 52274
rect 12798 52210 12850 52222
rect 32846 52210 32898 52222
rect 8990 52162 9042 52174
rect 8990 52098 9042 52110
rect 9998 52162 10050 52174
rect 9998 52098 10050 52110
rect 10334 52162 10386 52174
rect 11118 52162 11170 52174
rect 12350 52162 12402 52174
rect 10770 52110 10782 52162
rect 10834 52110 10846 52162
rect 11330 52110 11342 52162
rect 11394 52110 11406 52162
rect 11890 52110 11902 52162
rect 11954 52110 11966 52162
rect 10334 52098 10386 52110
rect 11118 52098 11170 52110
rect 12350 52098 12402 52110
rect 14590 52162 14642 52174
rect 14590 52098 14642 52110
rect 14814 52162 14866 52174
rect 14814 52098 14866 52110
rect 15598 52162 15650 52174
rect 15598 52098 15650 52110
rect 16270 52162 16322 52174
rect 27694 52162 27746 52174
rect 42590 52162 42642 52174
rect 20626 52110 20638 52162
rect 20690 52110 20702 52162
rect 27234 52110 27246 52162
rect 27298 52110 27310 52162
rect 29362 52110 29374 52162
rect 29426 52110 29438 52162
rect 33506 52110 33518 52162
rect 33570 52110 33582 52162
rect 38322 52110 38334 52162
rect 38386 52110 38398 52162
rect 40226 52110 40238 52162
rect 40290 52110 40302 52162
rect 41458 52110 41470 52162
rect 41522 52110 41534 52162
rect 41906 52110 41918 52162
rect 41970 52110 41982 52162
rect 43026 52110 43038 52162
rect 43090 52110 43102 52162
rect 16270 52098 16322 52110
rect 27694 52098 27746 52110
rect 42590 52098 42642 52110
rect 15150 52050 15202 52062
rect 41246 52050 41298 52062
rect 25218 51998 25230 52050
rect 25282 51998 25294 52050
rect 39218 51998 39230 52050
rect 39282 51998 39294 52050
rect 15150 51986 15202 51998
rect 41246 51986 41298 51998
rect 41358 52050 41410 52062
rect 41358 51986 41410 51998
rect 42254 52050 42306 52062
rect 42254 51986 42306 51998
rect 10110 51938 10162 51950
rect 10110 51874 10162 51886
rect 11902 51938 11954 51950
rect 11902 51874 11954 51886
rect 14702 51938 14754 51950
rect 14702 51874 14754 51886
rect 15710 51938 15762 51950
rect 15710 51874 15762 51886
rect 15822 51938 15874 51950
rect 15822 51874 15874 51886
rect 37102 51938 37154 51950
rect 37102 51874 37154 51886
rect 1344 51770 58576 51804
rect 1344 51718 19838 51770
rect 19890 51718 19942 51770
rect 19994 51718 20046 51770
rect 20098 51718 50558 51770
rect 50610 51718 50662 51770
rect 50714 51718 50766 51770
rect 50818 51718 58576 51770
rect 1344 51684 58576 51718
rect 12014 51602 12066 51614
rect 18174 51602 18226 51614
rect 16482 51550 16494 51602
rect 16546 51550 16558 51602
rect 17378 51550 17390 51602
rect 17442 51550 17454 51602
rect 12014 51538 12066 51550
rect 18174 51538 18226 51550
rect 18286 51602 18338 51614
rect 18286 51538 18338 51550
rect 18622 51602 18674 51614
rect 18622 51538 18674 51550
rect 40014 51602 40066 51614
rect 40014 51538 40066 51550
rect 41806 51602 41858 51614
rect 41806 51538 41858 51550
rect 42254 51602 42306 51614
rect 42254 51538 42306 51550
rect 2046 51490 2098 51502
rect 2046 51426 2098 51438
rect 10670 51490 10722 51502
rect 40238 51490 40290 51502
rect 10882 51438 10894 51490
rect 10946 51438 10958 51490
rect 13906 51438 13918 51490
rect 13970 51438 13982 51490
rect 21746 51438 21758 51490
rect 21810 51438 21822 51490
rect 10670 51426 10722 51438
rect 40238 51426 40290 51438
rect 41022 51490 41074 51502
rect 41234 51438 41246 51490
rect 41298 51438 41310 51490
rect 41022 51426 41074 51438
rect 7646 51378 7698 51390
rect 1810 51326 1822 51378
rect 1874 51326 1886 51378
rect 4386 51326 4398 51378
rect 4450 51326 4462 51378
rect 7646 51314 7698 51326
rect 11118 51378 11170 51390
rect 16830 51378 16882 51390
rect 11218 51326 11230 51378
rect 11282 51326 11294 51378
rect 13234 51326 13246 51378
rect 13298 51326 13310 51378
rect 11118 51314 11170 51326
rect 16830 51314 16882 51326
rect 17726 51378 17778 51390
rect 17726 51314 17778 51326
rect 18398 51378 18450 51390
rect 38446 51378 38498 51390
rect 21074 51326 21086 51378
rect 21138 51326 21150 51378
rect 25330 51326 25342 51378
rect 25394 51326 25406 51378
rect 18398 51314 18450 51326
rect 38446 51314 38498 51326
rect 38782 51378 38834 51390
rect 38994 51326 39006 51378
rect 39058 51326 39070 51378
rect 39554 51326 39566 51378
rect 39618 51326 39630 51378
rect 41794 51326 41806 51378
rect 41858 51326 41870 51378
rect 38782 51314 38834 51326
rect 2494 51266 2546 51278
rect 10782 51266 10834 51278
rect 38894 51266 38946 51278
rect 5058 51214 5070 51266
rect 5122 51214 5134 51266
rect 7186 51214 7198 51266
rect 7250 51214 7262 51266
rect 16034 51214 16046 51266
rect 16098 51214 16110 51266
rect 23874 51214 23886 51266
rect 23938 51214 23950 51266
rect 26114 51214 26126 51266
rect 26178 51214 26190 51266
rect 28242 51214 28254 51266
rect 28306 51214 28318 51266
rect 39890 51214 39902 51266
rect 39954 51214 39966 51266
rect 42130 51214 42142 51266
rect 42194 51214 42206 51266
rect 2494 51202 2546 51214
rect 10782 51202 10834 51214
rect 38894 51202 38946 51214
rect 39230 51154 39282 51166
rect 42478 51154 42530 51166
rect 41570 51102 41582 51154
rect 41634 51102 41646 51154
rect 39230 51090 39282 51102
rect 42478 51090 42530 51102
rect 1344 50986 58576 51020
rect 1344 50934 4478 50986
rect 4530 50934 4582 50986
rect 4634 50934 4686 50986
rect 4738 50934 35198 50986
rect 35250 50934 35302 50986
rect 35354 50934 35406 50986
rect 35458 50934 58576 50986
rect 1344 50900 58576 50934
rect 7310 50818 7362 50830
rect 7310 50754 7362 50766
rect 5070 50706 5122 50718
rect 1698 50654 1710 50706
rect 1762 50654 1774 50706
rect 3826 50654 3838 50706
rect 3890 50654 3902 50706
rect 5070 50642 5122 50654
rect 7086 50706 7138 50718
rect 7086 50642 7138 50654
rect 15934 50706 15986 50718
rect 15934 50642 15986 50654
rect 16494 50706 16546 50718
rect 16494 50642 16546 50654
rect 23662 50706 23714 50718
rect 23662 50642 23714 50654
rect 26462 50706 26514 50718
rect 26462 50642 26514 50654
rect 27358 50706 27410 50718
rect 27358 50642 27410 50654
rect 34526 50706 34578 50718
rect 40462 50706 40514 50718
rect 37874 50654 37886 50706
rect 37938 50654 37950 50706
rect 40002 50654 40014 50706
rect 40066 50654 40078 50706
rect 34526 50642 34578 50654
rect 40462 50642 40514 50654
rect 40910 50706 40962 50718
rect 42018 50654 42030 50706
rect 42082 50654 42094 50706
rect 44146 50654 44158 50706
rect 44210 50654 44222 50706
rect 40910 50642 40962 50654
rect 21870 50594 21922 50606
rect 4610 50542 4622 50594
rect 4674 50542 4686 50594
rect 21870 50530 21922 50542
rect 22094 50594 22146 50606
rect 22094 50530 22146 50542
rect 23774 50594 23826 50606
rect 23774 50530 23826 50542
rect 24446 50594 24498 50606
rect 24446 50530 24498 50542
rect 26238 50594 26290 50606
rect 26238 50530 26290 50542
rect 26686 50594 26738 50606
rect 26686 50530 26738 50542
rect 26798 50594 26850 50606
rect 26798 50530 26850 50542
rect 30382 50594 30434 50606
rect 35074 50542 35086 50594
rect 35138 50542 35150 50594
rect 37090 50542 37102 50594
rect 37154 50542 37166 50594
rect 41234 50542 41246 50594
rect 41298 50542 41310 50594
rect 30382 50530 30434 50542
rect 18174 50482 18226 50494
rect 23550 50482 23602 50494
rect 22418 50430 22430 50482
rect 22482 50430 22494 50482
rect 18174 50418 18226 50430
rect 23550 50418 23602 50430
rect 23998 50482 24050 50494
rect 24770 50430 24782 50482
rect 24834 50430 24846 50482
rect 23998 50418 24050 50430
rect 11902 50370 11954 50382
rect 7634 50318 7646 50370
rect 7698 50318 7710 50370
rect 11902 50306 11954 50318
rect 12574 50370 12626 50382
rect 12574 50306 12626 50318
rect 16046 50370 16098 50382
rect 16046 50306 16098 50318
rect 18286 50370 18338 50382
rect 18286 50306 18338 50318
rect 18510 50370 18562 50382
rect 32398 50370 32450 50382
rect 30706 50318 30718 50370
rect 30770 50318 30782 50370
rect 34850 50318 34862 50370
rect 34914 50318 34926 50370
rect 18510 50306 18562 50318
rect 32398 50306 32450 50318
rect 1344 50202 58576 50236
rect 1344 50150 19838 50202
rect 19890 50150 19942 50202
rect 19994 50150 20046 50202
rect 20098 50150 50558 50202
rect 50610 50150 50662 50202
rect 50714 50150 50766 50202
rect 50818 50150 58576 50202
rect 1344 50116 58576 50150
rect 5070 50034 5122 50046
rect 5070 49970 5122 49982
rect 7086 50034 7138 50046
rect 7086 49970 7138 49982
rect 11342 50034 11394 50046
rect 11342 49970 11394 49982
rect 12014 50034 12066 50046
rect 33070 50034 33122 50046
rect 13122 49982 13134 50034
rect 13186 49982 13198 50034
rect 12014 49970 12066 49982
rect 33070 49970 33122 49982
rect 41022 50034 41074 50046
rect 41022 49970 41074 49982
rect 7198 49922 7250 49934
rect 3826 49870 3838 49922
rect 3890 49870 3902 49922
rect 7198 49858 7250 49870
rect 7534 49922 7586 49934
rect 25230 49922 25282 49934
rect 17602 49870 17614 49922
rect 17666 49870 17678 49922
rect 7534 49858 7586 49870
rect 25230 49858 25282 49870
rect 27582 49922 27634 49934
rect 27582 49858 27634 49870
rect 8430 49810 8482 49822
rect 4610 49758 4622 49810
rect 4674 49758 4686 49810
rect 6514 49758 6526 49810
rect 6578 49758 6590 49810
rect 8430 49746 8482 49758
rect 8990 49810 9042 49822
rect 8990 49746 9042 49758
rect 10558 49810 10610 49822
rect 23102 49810 23154 49822
rect 33294 49810 33346 49822
rect 11554 49758 11566 49810
rect 11618 49758 11630 49810
rect 12226 49758 12238 49810
rect 12290 49758 12302 49810
rect 12898 49758 12910 49810
rect 12962 49758 12974 49810
rect 22642 49758 22654 49810
rect 22706 49758 22718 49810
rect 32162 49758 32174 49810
rect 32226 49758 32238 49810
rect 10558 49746 10610 49758
rect 23102 49746 23154 49758
rect 33294 49746 33346 49758
rect 33742 49810 33794 49822
rect 33742 49746 33794 49758
rect 34414 49810 34466 49822
rect 34414 49746 34466 49758
rect 34750 49810 34802 49822
rect 34750 49746 34802 49758
rect 35086 49810 35138 49822
rect 35086 49746 35138 49758
rect 8094 49698 8146 49710
rect 24110 49698 24162 49710
rect 33182 49698 33234 49710
rect 1698 49646 1710 49698
rect 1762 49646 1774 49698
rect 10098 49646 10110 49698
rect 10162 49646 10174 49698
rect 29250 49646 29262 49698
rect 29314 49646 29326 49698
rect 31378 49646 31390 49698
rect 31442 49646 31454 49698
rect 8094 49634 8146 49646
rect 24110 49634 24162 49646
rect 33182 49634 33234 49646
rect 34862 49698 34914 49710
rect 34862 49634 34914 49646
rect 35422 49698 35474 49710
rect 35422 49634 35474 49646
rect 6414 49586 6466 49598
rect 6414 49522 6466 49534
rect 11230 49586 11282 49598
rect 11230 49522 11282 49534
rect 11902 49586 11954 49598
rect 11902 49522 11954 49534
rect 25342 49586 25394 49598
rect 25342 49522 25394 49534
rect 27694 49586 27746 49598
rect 27694 49522 27746 49534
rect 1344 49418 58576 49452
rect 1344 49366 4478 49418
rect 4530 49366 4582 49418
rect 4634 49366 4686 49418
rect 4738 49366 35198 49418
rect 35250 49366 35302 49418
rect 35354 49366 35406 49418
rect 35458 49366 58576 49418
rect 1344 49332 58576 49366
rect 11118 49250 11170 49262
rect 18734 49250 18786 49262
rect 15810 49198 15822 49250
rect 15874 49198 15886 49250
rect 11118 49186 11170 49198
rect 18734 49186 18786 49198
rect 10222 49138 10274 49150
rect 11902 49138 11954 49150
rect 24558 49138 24610 49150
rect 32958 49138 33010 49150
rect 11330 49086 11342 49138
rect 11394 49086 11406 49138
rect 15474 49086 15486 49138
rect 15538 49086 15550 49138
rect 19058 49086 19070 49138
rect 19122 49086 19134 49138
rect 29586 49086 29598 49138
rect 29650 49086 29662 49138
rect 33506 49086 33518 49138
rect 33570 49086 33582 49138
rect 35634 49086 35646 49138
rect 35698 49086 35710 49138
rect 10222 49074 10274 49086
rect 11902 49074 11954 49086
rect 24558 49074 24610 49086
rect 32958 49074 33010 49086
rect 6526 49026 6578 49038
rect 22094 49026 22146 49038
rect 6962 48974 6974 49026
rect 7026 48974 7038 49026
rect 11442 48974 11454 49026
rect 11506 48974 11518 49026
rect 15362 48974 15374 49026
rect 15426 48974 15438 49026
rect 18162 48974 18174 49026
rect 18226 48974 18238 49026
rect 21858 48974 21870 49026
rect 21922 48974 21934 49026
rect 6526 48962 6578 48974
rect 22094 48962 22146 48974
rect 22206 49026 22258 49038
rect 22206 48962 22258 48974
rect 24670 49026 24722 49038
rect 25554 48974 25566 49026
rect 25618 48974 25630 49026
rect 27234 48974 27246 49026
rect 27298 48974 27310 49026
rect 32498 48974 32510 49026
rect 32562 48974 32574 49026
rect 36418 48974 36430 49026
rect 36482 48974 36494 49026
rect 24670 48962 24722 48974
rect 1710 48914 1762 48926
rect 1710 48850 1762 48862
rect 16382 48914 16434 48926
rect 16382 48850 16434 48862
rect 16494 48914 16546 48926
rect 16494 48850 16546 48862
rect 20414 48914 20466 48926
rect 20414 48850 20466 48862
rect 20526 48914 20578 48926
rect 20526 48850 20578 48862
rect 22542 48914 22594 48926
rect 22542 48850 22594 48862
rect 22878 48914 22930 48926
rect 22878 48850 22930 48862
rect 22990 48914 23042 48926
rect 26002 48862 26014 48914
rect 26066 48862 26078 48914
rect 27794 48862 27806 48914
rect 27858 48862 27870 48914
rect 31714 48862 31726 48914
rect 31778 48862 31790 48914
rect 22990 48850 23042 48862
rect 2046 48802 2098 48814
rect 2046 48738 2098 48750
rect 2494 48802 2546 48814
rect 2494 48738 2546 48750
rect 9662 48802 9714 48814
rect 9662 48738 9714 48750
rect 12462 48802 12514 48814
rect 12462 48738 12514 48750
rect 14478 48802 14530 48814
rect 14478 48738 14530 48750
rect 14926 48802 14978 48814
rect 14926 48738 14978 48750
rect 16158 48802 16210 48814
rect 18958 48802 19010 48814
rect 18386 48750 18398 48802
rect 18450 48750 18462 48802
rect 16158 48738 16210 48750
rect 18958 48738 19010 48750
rect 19630 48802 19682 48814
rect 19630 48738 19682 48750
rect 20190 48802 20242 48814
rect 20190 48738 20242 48750
rect 22430 48802 22482 48814
rect 22430 48738 22482 48750
rect 23214 48802 23266 48814
rect 37102 48802 37154 48814
rect 27122 48750 27134 48802
rect 27186 48750 27198 48802
rect 23214 48738 23266 48750
rect 37102 48738 37154 48750
rect 38894 48802 38946 48814
rect 38894 48738 38946 48750
rect 1344 48634 58576 48668
rect 1344 48582 19838 48634
rect 19890 48582 19942 48634
rect 19994 48582 20046 48634
rect 20098 48582 50558 48634
rect 50610 48582 50662 48634
rect 50714 48582 50766 48634
rect 50818 48582 58576 48634
rect 1344 48548 58576 48582
rect 3502 48466 3554 48478
rect 3502 48402 3554 48414
rect 16606 48466 16658 48478
rect 16606 48402 16658 48414
rect 22878 48466 22930 48478
rect 22878 48402 22930 48414
rect 30494 48466 30546 48478
rect 30494 48402 30546 48414
rect 31390 48466 31442 48478
rect 31390 48402 31442 48414
rect 39230 48466 39282 48478
rect 39230 48402 39282 48414
rect 7086 48354 7138 48366
rect 7086 48290 7138 48302
rect 7198 48354 7250 48366
rect 7198 48290 7250 48302
rect 10782 48354 10834 48366
rect 23438 48354 23490 48366
rect 19282 48302 19294 48354
rect 19346 48302 19358 48354
rect 19618 48302 19630 48354
rect 19682 48302 19694 48354
rect 21858 48302 21870 48354
rect 21922 48302 21934 48354
rect 10782 48290 10834 48302
rect 23438 48290 23490 48302
rect 23886 48354 23938 48366
rect 23886 48290 23938 48302
rect 23998 48354 24050 48366
rect 23998 48290 24050 48302
rect 26462 48354 26514 48366
rect 31502 48354 31554 48366
rect 27346 48302 27358 48354
rect 27410 48302 27422 48354
rect 29474 48302 29486 48354
rect 29538 48302 29550 48354
rect 30818 48302 30830 48354
rect 30882 48302 30894 48354
rect 26462 48290 26514 48302
rect 31502 48290 31554 48302
rect 31726 48354 31778 48366
rect 38546 48302 38558 48354
rect 38610 48302 38622 48354
rect 39554 48302 39566 48354
rect 39618 48302 39630 48354
rect 31726 48290 31778 48302
rect 6638 48242 6690 48254
rect 6638 48178 6690 48190
rect 9662 48242 9714 48254
rect 14142 48242 14194 48254
rect 10546 48190 10558 48242
rect 10610 48190 10622 48242
rect 11330 48190 11342 48242
rect 11394 48190 11406 48242
rect 11778 48190 11790 48242
rect 11842 48190 11854 48242
rect 9662 48178 9714 48190
rect 14142 48178 14194 48190
rect 15374 48242 15426 48254
rect 20078 48242 20130 48254
rect 22766 48242 22818 48254
rect 18162 48190 18174 48242
rect 18226 48190 18238 48242
rect 18610 48190 18622 48242
rect 18674 48190 18686 48242
rect 21634 48190 21646 48242
rect 21698 48190 21710 48242
rect 15374 48178 15426 48190
rect 20078 48178 20130 48190
rect 22766 48178 22818 48190
rect 23102 48242 23154 48254
rect 23102 48178 23154 48190
rect 23326 48242 23378 48254
rect 23326 48178 23378 48190
rect 23662 48242 23714 48254
rect 23662 48178 23714 48190
rect 24558 48242 24610 48254
rect 24558 48178 24610 48190
rect 26574 48242 26626 48254
rect 29822 48242 29874 48254
rect 27122 48190 27134 48242
rect 27186 48190 27198 48242
rect 29026 48190 29038 48242
rect 29090 48190 29102 48242
rect 26574 48178 26626 48190
rect 29822 48178 29874 48190
rect 31166 48242 31218 48254
rect 33618 48190 33630 48242
rect 33682 48190 33694 48242
rect 31166 48178 31218 48190
rect 4062 48130 4114 48142
rect 4062 48066 4114 48078
rect 6078 48130 6130 48142
rect 6078 48066 6130 48078
rect 10222 48130 10274 48142
rect 10222 48066 10274 48078
rect 14366 48130 14418 48142
rect 16158 48130 16210 48142
rect 15250 48078 15262 48130
rect 15314 48078 15326 48130
rect 14366 48066 14418 48078
rect 16158 48066 16210 48078
rect 17614 48130 17666 48142
rect 17614 48066 17666 48078
rect 18734 48130 18786 48142
rect 18734 48066 18786 48078
rect 20302 48130 20354 48142
rect 20302 48066 20354 48078
rect 22430 48130 22482 48142
rect 22430 48066 22482 48078
rect 32174 48130 32226 48142
rect 32174 48066 32226 48078
rect 33294 48130 33346 48142
rect 33294 48066 33346 48078
rect 7086 48018 7138 48030
rect 13470 48018 13522 48030
rect 11666 47966 11678 48018
rect 11730 47966 11742 48018
rect 7086 47954 7138 47966
rect 13470 47954 13522 47966
rect 13918 48018 13970 48030
rect 17502 48018 17554 48030
rect 15586 47966 15598 48018
rect 15650 47966 15662 48018
rect 16146 47966 16158 48018
rect 16210 48015 16222 48018
rect 16370 48015 16382 48018
rect 16210 47969 16382 48015
rect 16210 47966 16222 47969
rect 16370 47966 16382 47969
rect 16434 47966 16446 48018
rect 13918 47954 13970 47966
rect 17502 47954 17554 47966
rect 23998 48018 24050 48030
rect 23998 47954 24050 47966
rect 1344 47850 58576 47884
rect 1344 47798 4478 47850
rect 4530 47798 4582 47850
rect 4634 47798 4686 47850
rect 4738 47798 35198 47850
rect 35250 47798 35302 47850
rect 35354 47798 35406 47850
rect 35458 47798 58576 47850
rect 1344 47764 58576 47798
rect 3278 47682 3330 47694
rect 18510 47682 18562 47694
rect 16146 47630 16158 47682
rect 16210 47679 16222 47682
rect 16818 47679 16830 47682
rect 16210 47633 16830 47679
rect 16210 47630 16222 47633
rect 16818 47630 16830 47633
rect 16882 47630 16894 47682
rect 3278 47618 3330 47630
rect 18510 47618 18562 47630
rect 19294 47682 19346 47694
rect 19294 47618 19346 47630
rect 16830 47570 16882 47582
rect 2594 47518 2606 47570
rect 2658 47518 2670 47570
rect 7746 47518 7758 47570
rect 7810 47518 7822 47570
rect 16830 47506 16882 47518
rect 18174 47570 18226 47582
rect 18174 47506 18226 47518
rect 32062 47570 32114 47582
rect 32062 47506 32114 47518
rect 32846 47570 32898 47582
rect 32846 47506 32898 47518
rect 34302 47570 34354 47582
rect 34302 47506 34354 47518
rect 35758 47570 35810 47582
rect 35758 47506 35810 47518
rect 37774 47570 37826 47582
rect 39890 47518 39902 47570
rect 39954 47518 39966 47570
rect 37774 47506 37826 47518
rect 2158 47458 2210 47470
rect 2158 47394 2210 47406
rect 3950 47458 4002 47470
rect 7310 47458 7362 47470
rect 8766 47458 8818 47470
rect 6626 47406 6638 47458
rect 6690 47406 6702 47458
rect 8306 47406 8318 47458
rect 8370 47406 8382 47458
rect 3950 47394 4002 47406
rect 7310 47394 7362 47406
rect 8766 47394 8818 47406
rect 10782 47458 10834 47470
rect 10782 47394 10834 47406
rect 12798 47458 12850 47470
rect 12798 47394 12850 47406
rect 13582 47458 13634 47470
rect 13582 47394 13634 47406
rect 13806 47458 13858 47470
rect 13806 47394 13858 47406
rect 14030 47458 14082 47470
rect 15710 47458 15762 47470
rect 14802 47406 14814 47458
rect 14866 47406 14878 47458
rect 15362 47406 15374 47458
rect 15426 47406 15438 47458
rect 14030 47394 14082 47406
rect 15710 47394 15762 47406
rect 16046 47458 16098 47470
rect 16046 47394 16098 47406
rect 17166 47458 17218 47470
rect 17166 47394 17218 47406
rect 18286 47458 18338 47470
rect 19518 47458 19570 47470
rect 19170 47406 19182 47458
rect 19234 47406 19246 47458
rect 18286 47394 18338 47406
rect 19518 47394 19570 47406
rect 19742 47458 19794 47470
rect 33182 47458 33234 47470
rect 20066 47406 20078 47458
rect 20130 47406 20142 47458
rect 25890 47406 25902 47458
rect 25954 47406 25966 47458
rect 27346 47406 27358 47458
rect 27410 47406 27422 47458
rect 29362 47406 29374 47458
rect 29426 47406 29438 47458
rect 30930 47406 30942 47458
rect 30994 47406 31006 47458
rect 31266 47406 31278 47458
rect 31330 47406 31342 47458
rect 19742 47394 19794 47406
rect 33182 47394 33234 47406
rect 33742 47458 33794 47470
rect 33742 47394 33794 47406
rect 34190 47458 34242 47470
rect 34190 47394 34242 47406
rect 34974 47458 35026 47470
rect 34974 47394 35026 47406
rect 35310 47458 35362 47470
rect 35310 47394 35362 47406
rect 38110 47458 38162 47470
rect 38110 47394 38162 47406
rect 39006 47458 39058 47470
rect 42690 47406 42702 47458
rect 42754 47406 42766 47458
rect 39006 47394 39058 47406
rect 3054 47346 3106 47358
rect 3054 47282 3106 47294
rect 4510 47346 4562 47358
rect 4510 47282 4562 47294
rect 6190 47346 6242 47358
rect 12238 47346 12290 47358
rect 9202 47294 9214 47346
rect 9266 47294 9278 47346
rect 6190 47282 6242 47294
rect 12238 47282 12290 47294
rect 17278 47346 17330 47358
rect 17278 47282 17330 47294
rect 18958 47346 19010 47358
rect 34750 47346 34802 47358
rect 26002 47294 26014 47346
rect 26066 47294 26078 47346
rect 28130 47294 28142 47346
rect 28194 47294 28206 47346
rect 29138 47294 29150 47346
rect 29202 47294 29214 47346
rect 33506 47294 33518 47346
rect 33570 47294 33582 47346
rect 42018 47294 42030 47346
rect 42082 47294 42094 47346
rect 18958 47282 19010 47294
rect 34750 47282 34802 47294
rect 14478 47234 14530 47246
rect 3602 47182 3614 47234
rect 3666 47182 3678 47234
rect 12674 47182 12686 47234
rect 12738 47182 12750 47234
rect 14478 47170 14530 47182
rect 16382 47234 16434 47246
rect 16382 47170 16434 47182
rect 17502 47234 17554 47246
rect 17502 47170 17554 47182
rect 18174 47234 18226 47246
rect 18174 47170 18226 47182
rect 20302 47234 20354 47246
rect 20302 47170 20354 47182
rect 20414 47234 20466 47246
rect 20414 47170 20466 47182
rect 24670 47234 24722 47246
rect 34414 47234 34466 47246
rect 26898 47182 26910 47234
rect 26962 47182 26974 47234
rect 24670 47170 24722 47182
rect 34414 47170 34466 47182
rect 35198 47234 35250 47246
rect 39118 47234 39170 47246
rect 38434 47182 38446 47234
rect 38498 47182 38510 47234
rect 35198 47170 35250 47182
rect 39118 47170 39170 47182
rect 39230 47234 39282 47246
rect 39230 47170 39282 47182
rect 39454 47234 39506 47246
rect 39454 47170 39506 47182
rect 1344 47066 58576 47100
rect 1344 47014 19838 47066
rect 19890 47014 19942 47066
rect 19994 47014 20046 47066
rect 20098 47014 50558 47066
rect 50610 47014 50662 47066
rect 50714 47014 50766 47066
rect 50818 47014 58576 47066
rect 1344 46980 58576 47014
rect 2494 46898 2546 46910
rect 16158 46898 16210 46910
rect 13346 46846 13358 46898
rect 13410 46846 13422 46898
rect 2494 46834 2546 46846
rect 16158 46834 16210 46846
rect 33406 46898 33458 46910
rect 33406 46834 33458 46846
rect 38894 46898 38946 46910
rect 38894 46834 38946 46846
rect 40014 46898 40066 46910
rect 40014 46834 40066 46846
rect 40350 46898 40402 46910
rect 40350 46834 40402 46846
rect 41246 46898 41298 46910
rect 41246 46834 41298 46846
rect 1710 46786 1762 46798
rect 1710 46722 1762 46734
rect 2046 46786 2098 46798
rect 2046 46722 2098 46734
rect 2942 46786 2994 46798
rect 6414 46786 6466 46798
rect 3714 46734 3726 46786
rect 3778 46734 3790 46786
rect 4834 46734 4846 46786
rect 4898 46734 4910 46786
rect 2942 46722 2994 46734
rect 6414 46722 6466 46734
rect 7870 46786 7922 46798
rect 13134 46786 13186 46798
rect 10322 46734 10334 46786
rect 10386 46734 10398 46786
rect 11330 46734 11342 46786
rect 11394 46734 11406 46786
rect 7870 46722 7922 46734
rect 13134 46722 13186 46734
rect 19966 46786 20018 46798
rect 33630 46786 33682 46798
rect 40910 46786 40962 46798
rect 27906 46734 27918 46786
rect 27970 46734 27982 46786
rect 36642 46734 36654 46786
rect 36706 46734 36718 46786
rect 39442 46734 39454 46786
rect 39506 46734 39518 46786
rect 19966 46722 20018 46734
rect 33630 46722 33682 46734
rect 40910 46722 40962 46734
rect 41134 46786 41186 46798
rect 41134 46722 41186 46734
rect 41470 46786 41522 46798
rect 41470 46722 41522 46734
rect 4510 46674 4562 46686
rect 7310 46674 7362 46686
rect 15038 46674 15090 46686
rect 32622 46674 32674 46686
rect 3938 46622 3950 46674
rect 4002 46622 4014 46674
rect 6962 46622 6974 46674
rect 7026 46622 7038 46674
rect 10434 46622 10446 46674
rect 10498 46622 10510 46674
rect 11442 46622 11454 46674
rect 11506 46622 11518 46674
rect 13570 46622 13582 46674
rect 13634 46622 13646 46674
rect 14130 46622 14142 46674
rect 14194 46622 14206 46674
rect 14690 46622 14702 46674
rect 14754 46622 14766 46674
rect 20290 46622 20302 46674
rect 20354 46622 20366 46674
rect 25218 46622 25230 46674
rect 25282 46622 25294 46674
rect 4510 46610 4562 46622
rect 7310 46610 7362 46622
rect 15038 46610 15090 46622
rect 32622 46610 32674 46622
rect 33070 46674 33122 46686
rect 33070 46610 33122 46622
rect 33294 46674 33346 46686
rect 39118 46674 39170 46686
rect 37314 46622 37326 46674
rect 37378 46622 37390 46674
rect 33294 46610 33346 46622
rect 39118 46610 39170 46622
rect 15710 46562 15762 46574
rect 3826 46510 3838 46562
rect 3890 46510 3902 46562
rect 5954 46510 5966 46562
rect 6018 46510 6030 46562
rect 15710 46498 15762 46510
rect 22766 46562 22818 46574
rect 22766 46498 22818 46510
rect 24334 46562 24386 46574
rect 24334 46498 24386 46510
rect 24782 46562 24834 46574
rect 34514 46510 34526 46562
rect 34578 46510 34590 46562
rect 24782 46498 24834 46510
rect 3054 46450 3106 46462
rect 20302 46450 20354 46462
rect 15026 46398 15038 46450
rect 15090 46398 15102 46450
rect 3054 46386 3106 46398
rect 20302 46386 20354 46398
rect 1344 46282 58576 46316
rect 1344 46230 4478 46282
rect 4530 46230 4582 46282
rect 4634 46230 4686 46282
rect 4738 46230 35198 46282
rect 35250 46230 35302 46282
rect 35354 46230 35406 46282
rect 35458 46230 58576 46282
rect 1344 46196 58576 46230
rect 14690 46062 14702 46114
rect 14754 46111 14766 46114
rect 15026 46111 15038 46114
rect 14754 46065 15038 46111
rect 14754 46062 14766 46065
rect 15026 46062 15038 46065
rect 15090 46062 15102 46114
rect 9886 46002 9938 46014
rect 7298 45950 7310 46002
rect 7362 45950 7374 46002
rect 9886 45938 9938 45950
rect 14478 46002 14530 46014
rect 14478 45938 14530 45950
rect 15038 46002 15090 46014
rect 15038 45938 15090 45950
rect 22206 46002 22258 46014
rect 22206 45938 22258 45950
rect 22654 46002 22706 46014
rect 32062 46002 32114 46014
rect 27794 45950 27806 46002
rect 27858 45950 27870 46002
rect 22654 45938 22706 45950
rect 32062 45938 32114 45950
rect 32846 46002 32898 46014
rect 32846 45938 32898 45950
rect 33742 46002 33794 46014
rect 33742 45938 33794 45950
rect 34750 46002 34802 46014
rect 34750 45938 34802 45950
rect 41022 46002 41074 46014
rect 41022 45938 41074 45950
rect 3950 45890 4002 45902
rect 8654 45890 8706 45902
rect 12126 45890 12178 45902
rect 6850 45838 6862 45890
rect 6914 45838 6926 45890
rect 7634 45838 7646 45890
rect 7698 45838 7710 45890
rect 10322 45838 10334 45890
rect 10386 45838 10398 45890
rect 3950 45826 4002 45838
rect 8654 45826 8706 45838
rect 12126 45826 12178 45838
rect 13918 45890 13970 45902
rect 13918 45826 13970 45838
rect 16046 45890 16098 45902
rect 19966 45890 20018 45902
rect 16482 45838 16494 45890
rect 16546 45838 16558 45890
rect 16706 45838 16718 45890
rect 16770 45838 16782 45890
rect 16046 45826 16098 45838
rect 19966 45826 20018 45838
rect 20078 45890 20130 45902
rect 20078 45826 20130 45838
rect 21646 45890 21698 45902
rect 21646 45826 21698 45838
rect 21982 45890 22034 45902
rect 21982 45826 22034 45838
rect 24446 45890 24498 45902
rect 32734 45890 32786 45902
rect 24770 45838 24782 45890
rect 24834 45838 24846 45890
rect 26786 45838 26798 45890
rect 26850 45838 26862 45890
rect 29362 45838 29374 45890
rect 29426 45838 29438 45890
rect 31826 45838 31838 45890
rect 31890 45838 31902 45890
rect 24446 45826 24498 45838
rect 32734 45826 32786 45838
rect 32958 45890 33010 45902
rect 32958 45826 33010 45838
rect 33406 45890 33458 45902
rect 33406 45826 33458 45838
rect 34190 45890 34242 45902
rect 34190 45826 34242 45838
rect 34638 45890 34690 45902
rect 34638 45826 34690 45838
rect 34862 45890 34914 45902
rect 34862 45826 34914 45838
rect 38558 45890 38610 45902
rect 38558 45826 38610 45838
rect 38670 45890 38722 45902
rect 38670 45826 38722 45838
rect 41582 45890 41634 45902
rect 41582 45826 41634 45838
rect 41918 45890 41970 45902
rect 41918 45826 41970 45838
rect 1710 45778 1762 45790
rect 1710 45714 1762 45726
rect 4510 45778 4562 45790
rect 4510 45714 4562 45726
rect 6526 45778 6578 45790
rect 6526 45714 6578 45726
rect 9326 45778 9378 45790
rect 9326 45714 9378 45726
rect 10894 45778 10946 45790
rect 10894 45714 10946 45726
rect 16270 45778 16322 45790
rect 16270 45714 16322 45726
rect 17838 45778 17890 45790
rect 24558 45778 24610 45790
rect 27358 45778 27410 45790
rect 41358 45778 41410 45790
rect 23650 45726 23662 45778
rect 23714 45726 23726 45778
rect 24210 45726 24222 45778
rect 24274 45726 24286 45778
rect 24882 45726 24894 45778
rect 24946 45726 24958 45778
rect 29474 45726 29486 45778
rect 29538 45726 29550 45778
rect 31714 45726 31726 45778
rect 31778 45726 31790 45778
rect 17838 45714 17890 45726
rect 24558 45714 24610 45726
rect 27358 45714 27410 45726
rect 41358 45714 41410 45726
rect 2046 45666 2098 45678
rect 2046 45602 2098 45614
rect 2494 45666 2546 45678
rect 2494 45602 2546 45614
rect 6638 45666 6690 45678
rect 6638 45602 6690 45614
rect 8094 45666 8146 45678
rect 8094 45602 8146 45614
rect 10446 45666 10498 45678
rect 10446 45602 10498 45614
rect 16158 45666 16210 45678
rect 16158 45602 16210 45614
rect 17390 45666 17442 45678
rect 17390 45602 17442 45614
rect 19742 45666 19794 45678
rect 19742 45602 19794 45614
rect 20638 45666 20690 45678
rect 20638 45602 20690 45614
rect 21422 45666 21474 45678
rect 21422 45602 21474 45614
rect 21534 45666 21586 45678
rect 23102 45666 23154 45678
rect 22418 45614 22430 45666
rect 22482 45614 22494 45666
rect 21534 45602 21586 45614
rect 23102 45602 23154 45614
rect 41806 45666 41858 45678
rect 41806 45602 41858 45614
rect 1344 45498 58576 45532
rect 1344 45446 19838 45498
rect 19890 45446 19942 45498
rect 19994 45446 20046 45498
rect 20098 45446 50558 45498
rect 50610 45446 50662 45498
rect 50714 45446 50766 45498
rect 50818 45446 58576 45498
rect 1344 45412 58576 45446
rect 2606 45330 2658 45342
rect 2606 45266 2658 45278
rect 3166 45330 3218 45342
rect 3166 45266 3218 45278
rect 8206 45330 8258 45342
rect 21422 45330 21474 45342
rect 19058 45278 19070 45330
rect 19122 45278 19134 45330
rect 8206 45266 8258 45278
rect 21422 45266 21474 45278
rect 22654 45330 22706 45342
rect 25678 45330 25730 45342
rect 32510 45330 32562 45342
rect 23426 45278 23438 45330
rect 23490 45278 23502 45330
rect 27570 45278 27582 45330
rect 27634 45278 27646 45330
rect 22654 45266 22706 45278
rect 25678 45266 25730 45278
rect 32510 45266 32562 45278
rect 40238 45330 40290 45342
rect 40238 45266 40290 45278
rect 7982 45218 8034 45230
rect 7982 45154 8034 45166
rect 10222 45218 10274 45230
rect 21646 45218 21698 45230
rect 19394 45166 19406 45218
rect 19458 45166 19470 45218
rect 19618 45166 19630 45218
rect 19682 45166 19694 45218
rect 10222 45154 10274 45166
rect 21646 45154 21698 45166
rect 22542 45218 22594 45230
rect 22542 45154 22594 45166
rect 25902 45218 25954 45230
rect 28702 45218 28754 45230
rect 26226 45166 26238 45218
rect 26290 45166 26302 45218
rect 25902 45154 25954 45166
rect 28702 45154 28754 45166
rect 33182 45218 33234 45230
rect 33182 45154 33234 45166
rect 33406 45218 33458 45230
rect 42354 45166 42366 45218
rect 42418 45166 42430 45218
rect 33406 45154 33458 45166
rect 2494 45106 2546 45118
rect 2494 45042 2546 45054
rect 2830 45106 2882 45118
rect 2830 45042 2882 45054
rect 3054 45106 3106 45118
rect 6862 45106 6914 45118
rect 7758 45106 7810 45118
rect 4162 45054 4174 45106
rect 4226 45054 4238 45106
rect 6962 45054 6974 45106
rect 7026 45054 7038 45106
rect 3054 45042 3106 45054
rect 6862 45042 6914 45054
rect 7758 45042 7810 45054
rect 11118 45106 11170 45118
rect 11118 45042 11170 45054
rect 11454 45106 11506 45118
rect 11454 45042 11506 45054
rect 13806 45106 13858 45118
rect 20750 45106 20802 45118
rect 22318 45106 22370 45118
rect 19954 45054 19966 45106
rect 20018 45054 20030 45106
rect 21858 45054 21870 45106
rect 21922 45054 21934 45106
rect 13806 45042 13858 45054
rect 20750 45042 20802 45054
rect 22318 45042 22370 45054
rect 22878 45106 22930 45118
rect 22878 45042 22930 45054
rect 25566 45106 25618 45118
rect 39678 45106 39730 45118
rect 26114 45054 26126 45106
rect 26178 45054 26190 45106
rect 29922 45054 29934 45106
rect 29986 45054 29998 45106
rect 33842 45054 33854 45106
rect 33906 45054 33918 45106
rect 25566 45042 25618 45054
rect 39678 45042 39730 45054
rect 40126 45106 40178 45118
rect 40126 45042 40178 45054
rect 40350 45106 40402 45118
rect 41570 45054 41582 45106
rect 41634 45054 41646 45106
rect 40350 45042 40402 45054
rect 11566 44994 11618 45006
rect 3826 44942 3838 44994
rect 3890 44942 3902 44994
rect 6738 44942 6750 44994
rect 6802 44942 6814 44994
rect 8194 44942 8206 44994
rect 8258 44942 8270 44994
rect 11566 44930 11618 44942
rect 14366 44994 14418 45006
rect 14366 44930 14418 44942
rect 18622 44994 18674 45006
rect 18622 44930 18674 44942
rect 20302 44994 20354 45006
rect 20302 44930 20354 44942
rect 24334 44994 24386 45006
rect 24334 44930 24386 44942
rect 24670 44994 24722 45006
rect 36978 44942 36990 44994
rect 37042 44942 37054 44994
rect 44482 44942 44494 44994
rect 44546 44942 44558 44994
rect 24670 44930 24722 44942
rect 3166 44882 3218 44894
rect 3166 44818 3218 44830
rect 20526 44882 20578 44894
rect 20526 44818 20578 44830
rect 20974 44882 21026 44894
rect 20974 44818 21026 44830
rect 22094 44882 22146 44894
rect 22094 44818 22146 44830
rect 23102 44882 23154 44894
rect 23102 44818 23154 44830
rect 33518 44882 33570 44894
rect 33518 44818 33570 44830
rect 1344 44714 58576 44748
rect 1344 44662 4478 44714
rect 4530 44662 4582 44714
rect 4634 44662 4686 44714
rect 4738 44662 35198 44714
rect 35250 44662 35302 44714
rect 35354 44662 35406 44714
rect 35458 44662 58576 44714
rect 1344 44628 58576 44662
rect 25790 44546 25842 44558
rect 22082 44494 22094 44546
rect 22146 44494 22158 44546
rect 25790 44482 25842 44494
rect 27134 44546 27186 44558
rect 34402 44494 34414 44546
rect 34466 44494 34478 44546
rect 27134 44482 27186 44494
rect 13806 44434 13858 44446
rect 8530 44382 8542 44434
rect 8594 44382 8606 44434
rect 13806 44370 13858 44382
rect 14814 44434 14866 44446
rect 14814 44370 14866 44382
rect 16158 44434 16210 44446
rect 26126 44434 26178 44446
rect 35422 44434 35474 44446
rect 23426 44382 23438 44434
rect 23490 44382 23502 44434
rect 24658 44382 24670 44434
rect 24722 44382 24734 44434
rect 28466 44382 28478 44434
rect 28530 44382 28542 44434
rect 29362 44382 29374 44434
rect 29426 44382 29438 44434
rect 16158 44370 16210 44382
rect 26126 44370 26178 44382
rect 35422 44370 35474 44382
rect 37550 44434 37602 44446
rect 37550 44370 37602 44382
rect 38558 44434 38610 44446
rect 38558 44370 38610 44382
rect 10222 44322 10274 44334
rect 14254 44322 14306 44334
rect 15710 44322 15762 44334
rect 6850 44270 6862 44322
rect 6914 44270 6926 44322
rect 10434 44270 10446 44322
rect 10498 44270 10510 44322
rect 10994 44270 11006 44322
rect 11058 44270 11070 44322
rect 11218 44270 11230 44322
rect 11282 44270 11294 44322
rect 11442 44270 11454 44322
rect 11506 44270 11518 44322
rect 15250 44270 15262 44322
rect 15314 44270 15326 44322
rect 10222 44258 10274 44270
rect 14254 44258 14306 44270
rect 15710 44258 15762 44270
rect 16382 44322 16434 44334
rect 16382 44258 16434 44270
rect 16606 44322 16658 44334
rect 16606 44258 16658 44270
rect 16830 44322 16882 44334
rect 21646 44322 21698 44334
rect 17490 44270 17502 44322
rect 17554 44270 17566 44322
rect 20738 44270 20750 44322
rect 20802 44270 20814 44322
rect 21298 44270 21310 44322
rect 21362 44270 21374 44322
rect 16830 44258 16882 44270
rect 21646 44258 21698 44270
rect 22990 44322 23042 44334
rect 26350 44322 26402 44334
rect 29598 44322 29650 44334
rect 39006 44322 39058 44334
rect 24434 44270 24446 44322
rect 24498 44270 24510 44322
rect 26674 44270 26686 44322
rect 26738 44270 26750 44322
rect 30818 44270 30830 44322
rect 30882 44270 30894 44322
rect 33282 44270 33294 44322
rect 33346 44270 33358 44322
rect 34178 44270 34190 44322
rect 34242 44270 34254 44322
rect 34738 44270 34750 44322
rect 34802 44270 34814 44322
rect 22990 44258 23042 44270
rect 26350 44258 26402 44270
rect 29598 44258 29650 44270
rect 39006 44258 39058 44270
rect 39118 44322 39170 44334
rect 39118 44258 39170 44270
rect 39566 44322 39618 44334
rect 39566 44258 39618 44270
rect 8094 44210 8146 44222
rect 5730 44158 5742 44210
rect 5794 44158 5806 44210
rect 8094 44146 8146 44158
rect 10558 44210 10610 44222
rect 10558 44146 10610 44158
rect 17390 44210 17442 44222
rect 21534 44210 21586 44222
rect 19170 44158 19182 44210
rect 19234 44158 19246 44210
rect 19842 44158 19854 44210
rect 19906 44158 19918 44210
rect 17390 44146 17442 44158
rect 21534 44146 21586 44158
rect 22654 44210 22706 44222
rect 26462 44210 26514 44222
rect 24210 44158 24222 44210
rect 24274 44158 24286 44210
rect 22654 44146 22706 44158
rect 26462 44146 26514 44158
rect 29934 44210 29986 44222
rect 34974 44210 35026 44222
rect 30594 44158 30606 44210
rect 30658 44158 30670 44210
rect 32946 44158 32958 44210
rect 33010 44158 33022 44210
rect 29934 44146 29986 44158
rect 34974 44146 35026 44158
rect 37438 44210 37490 44222
rect 37438 44146 37490 44158
rect 12238 44098 12290 44110
rect 12238 44034 12290 44046
rect 17278 44098 17330 44110
rect 17278 44034 17330 44046
rect 25006 44098 25058 44110
rect 25006 44034 25058 44046
rect 27470 44098 27522 44110
rect 27470 44034 27522 44046
rect 27806 44098 27858 44110
rect 39342 44098 39394 44110
rect 32610 44046 32622 44098
rect 32674 44046 32686 44098
rect 34626 44046 34638 44098
rect 34690 44046 34702 44098
rect 27806 44034 27858 44046
rect 39342 44034 39394 44046
rect 1344 43930 58576 43964
rect 1344 43878 19838 43930
rect 19890 43878 19942 43930
rect 19994 43878 20046 43930
rect 20098 43878 50558 43930
rect 50610 43878 50662 43930
rect 50714 43878 50766 43930
rect 50818 43878 58576 43930
rect 1344 43844 58576 43878
rect 7198 43762 7250 43774
rect 7198 43698 7250 43710
rect 13246 43762 13298 43774
rect 13246 43698 13298 43710
rect 17502 43762 17554 43774
rect 22306 43710 22318 43762
rect 22370 43710 22382 43762
rect 23762 43710 23774 43762
rect 23826 43710 23838 43762
rect 28242 43710 28254 43762
rect 28306 43710 28318 43762
rect 17502 43698 17554 43710
rect 2270 43650 2322 43662
rect 2270 43586 2322 43598
rect 2718 43650 2770 43662
rect 2718 43586 2770 43598
rect 5294 43650 5346 43662
rect 5294 43586 5346 43598
rect 6526 43650 6578 43662
rect 6526 43586 6578 43598
rect 7758 43650 7810 43662
rect 7758 43586 7810 43598
rect 11006 43650 11058 43662
rect 11006 43586 11058 43598
rect 13134 43650 13186 43662
rect 13134 43586 13186 43598
rect 17390 43650 17442 43662
rect 17390 43586 17442 43598
rect 17614 43650 17666 43662
rect 21758 43650 21810 43662
rect 18722 43598 18734 43650
rect 18786 43598 18798 43650
rect 17614 43586 17666 43598
rect 21758 43586 21810 43598
rect 24558 43650 24610 43662
rect 26238 43650 26290 43662
rect 29150 43650 29202 43662
rect 25330 43598 25342 43650
rect 25394 43598 25406 43650
rect 26562 43598 26574 43650
rect 26626 43598 26638 43650
rect 24558 43586 24610 43598
rect 26238 43586 26290 43598
rect 29150 43586 29202 43598
rect 31502 43650 31554 43662
rect 31502 43586 31554 43598
rect 31726 43650 31778 43662
rect 32622 43650 32674 43662
rect 32050 43598 32062 43650
rect 32114 43598 32126 43650
rect 31726 43586 31778 43598
rect 32622 43586 32674 43598
rect 33070 43650 33122 43662
rect 41246 43650 41298 43662
rect 33394 43598 33406 43650
rect 33458 43598 33470 43650
rect 34626 43598 34638 43650
rect 34690 43598 34702 43650
rect 39330 43598 39342 43650
rect 39394 43598 39406 43650
rect 33070 43586 33122 43598
rect 41246 43586 41298 43598
rect 2494 43538 2546 43550
rect 3502 43538 3554 43550
rect 10110 43538 10162 43550
rect 13918 43538 13970 43550
rect 23438 43538 23490 43550
rect 2930 43486 2942 43538
rect 2994 43486 3006 43538
rect 4834 43486 4846 43538
rect 4898 43486 4910 43538
rect 6850 43486 6862 43538
rect 6914 43486 6926 43538
rect 12786 43486 12798 43538
rect 12850 43486 12862 43538
rect 13458 43486 13470 43538
rect 13522 43486 13534 43538
rect 17826 43486 17838 43538
rect 17890 43486 17902 43538
rect 18162 43486 18174 43538
rect 18226 43486 18238 43538
rect 18610 43486 18622 43538
rect 18674 43486 18686 43538
rect 20626 43486 20638 43538
rect 20690 43486 20702 43538
rect 2494 43474 2546 43486
rect 3502 43474 3554 43486
rect 10110 43474 10162 43486
rect 13918 43474 13970 43486
rect 23438 43474 23490 43486
rect 24222 43538 24274 43550
rect 24222 43474 24274 43486
rect 25566 43538 25618 43550
rect 41134 43538 41186 43550
rect 25778 43486 25790 43538
rect 25842 43486 25854 43538
rect 28130 43486 28142 43538
rect 28194 43486 28206 43538
rect 28578 43486 28590 43538
rect 28642 43486 28654 43538
rect 33954 43486 33966 43538
rect 34018 43486 34030 43538
rect 40002 43486 40014 43538
rect 40066 43486 40078 43538
rect 25566 43474 25618 43486
rect 41134 43474 41186 43486
rect 41358 43538 41410 43550
rect 41682 43486 41694 43538
rect 41746 43486 41758 43538
rect 41358 43474 41410 43486
rect 1822 43426 1874 43438
rect 4062 43426 4114 43438
rect 5854 43426 5906 43438
rect 2818 43374 2830 43426
rect 2882 43374 2894 43426
rect 4498 43374 4510 43426
rect 4562 43374 4574 43426
rect 1822 43362 1874 43374
rect 4062 43362 4114 43374
rect 5854 43362 5906 43374
rect 9998 43426 10050 43438
rect 12462 43426 12514 43438
rect 11330 43374 11342 43426
rect 11394 43374 11406 43426
rect 9998 43362 10050 43374
rect 12462 43362 12514 43374
rect 14478 43426 14530 43438
rect 14478 43362 14530 43374
rect 23102 43426 23154 43438
rect 23102 43362 23154 43374
rect 25230 43426 25282 43438
rect 36754 43374 36766 43426
rect 36818 43374 36830 43426
rect 37202 43374 37214 43426
rect 37266 43374 37278 43426
rect 25230 43362 25282 43374
rect 6862 43314 6914 43326
rect 6862 43250 6914 43262
rect 9662 43314 9714 43326
rect 9662 43250 9714 43262
rect 9774 43314 9826 43326
rect 24670 43314 24722 43326
rect 11442 43262 11454 43314
rect 11506 43262 11518 43314
rect 9774 43250 9826 43262
rect 24670 43250 24722 43262
rect 1344 43146 58576 43180
rect 1344 43094 4478 43146
rect 4530 43094 4582 43146
rect 4634 43094 4686 43146
rect 4738 43094 35198 43146
rect 35250 43094 35302 43146
rect 35354 43094 35406 43146
rect 35458 43094 58576 43146
rect 1344 43060 58576 43094
rect 23998 42978 24050 42990
rect 8306 42926 8318 42978
rect 8370 42926 8382 42978
rect 22642 42926 22654 42978
rect 22706 42975 22718 42978
rect 23426 42975 23438 42978
rect 22706 42929 23438 42975
rect 22706 42926 22718 42929
rect 23426 42926 23438 42929
rect 23490 42926 23502 42978
rect 24994 42926 25006 42978
rect 25058 42926 25070 42978
rect 30034 42926 30046 42978
rect 30098 42926 30110 42978
rect 23998 42914 24050 42926
rect 23662 42866 23714 42878
rect 7970 42814 7982 42866
rect 8034 42814 8046 42866
rect 13906 42814 13918 42866
rect 13970 42814 13982 42866
rect 21746 42814 21758 42866
rect 21810 42814 21822 42866
rect 23662 42802 23714 42814
rect 38670 42866 38722 42878
rect 38670 42802 38722 42814
rect 39118 42866 39170 42878
rect 44034 42814 44046 42866
rect 44098 42814 44110 42866
rect 39118 42802 39170 42814
rect 8206 42754 8258 42766
rect 13470 42754 13522 42766
rect 1810 42702 1822 42754
rect 1874 42702 1886 42754
rect 7858 42702 7870 42754
rect 7922 42702 7934 42754
rect 8754 42702 8766 42754
rect 8818 42702 8830 42754
rect 10770 42702 10782 42754
rect 10834 42702 10846 42754
rect 8206 42690 8258 42702
rect 13470 42690 13522 42702
rect 17614 42754 17666 42766
rect 24446 42754 24498 42766
rect 18050 42702 18062 42754
rect 18114 42702 18126 42754
rect 17614 42690 17666 42702
rect 24446 42690 24498 42702
rect 24670 42754 24722 42766
rect 24670 42690 24722 42702
rect 25566 42754 25618 42766
rect 30270 42754 30322 42766
rect 38558 42754 38610 42766
rect 27794 42702 27806 42754
rect 27858 42702 27870 42754
rect 29362 42702 29374 42754
rect 29426 42702 29438 42754
rect 29922 42702 29934 42754
rect 29986 42702 29998 42754
rect 31042 42702 31054 42754
rect 31106 42702 31118 42754
rect 33506 42702 33518 42754
rect 33570 42702 33582 42754
rect 25566 42690 25618 42702
rect 30270 42690 30322 42702
rect 38558 42690 38610 42702
rect 39230 42754 39282 42766
rect 39230 42690 39282 42702
rect 40126 42754 40178 42766
rect 40126 42690 40178 42702
rect 40798 42754 40850 42766
rect 41122 42702 41134 42754
rect 41186 42702 41198 42754
rect 40798 42690 40850 42702
rect 2046 42642 2098 42654
rect 2046 42578 2098 42590
rect 2718 42642 2770 42654
rect 2718 42578 2770 42590
rect 2830 42642 2882 42654
rect 11902 42642 11954 42654
rect 8866 42590 8878 42642
rect 8930 42590 8942 42642
rect 2830 42578 2882 42590
rect 11902 42578 11954 42590
rect 23886 42642 23938 42654
rect 39006 42642 39058 42654
rect 25442 42590 25454 42642
rect 25506 42590 25518 42642
rect 27346 42590 27358 42642
rect 27410 42590 27422 42642
rect 30818 42590 30830 42642
rect 30882 42590 30894 42642
rect 32946 42590 32958 42642
rect 33010 42590 33022 42642
rect 23886 42578 23938 42590
rect 39006 42578 39058 42590
rect 39454 42642 39506 42654
rect 39454 42578 39506 42590
rect 40574 42642 40626 42654
rect 41906 42590 41918 42642
rect 41970 42590 41982 42642
rect 40574 42578 40626 42590
rect 3054 42530 3106 42542
rect 20750 42530 20802 42542
rect 10322 42478 10334 42530
rect 10386 42478 10398 42530
rect 3054 42466 3106 42478
rect 20750 42466 20802 42478
rect 21310 42530 21362 42542
rect 21310 42466 21362 42478
rect 22654 42530 22706 42542
rect 22654 42466 22706 42478
rect 23214 42530 23266 42542
rect 23214 42466 23266 42478
rect 23998 42530 24050 42542
rect 23998 42466 24050 42478
rect 28366 42530 28418 42542
rect 34638 42530 34690 42542
rect 32834 42478 32846 42530
rect 32898 42478 32910 42530
rect 28366 42466 28418 42478
rect 34638 42466 34690 42478
rect 40462 42530 40514 42542
rect 40462 42466 40514 42478
rect 1344 42362 58576 42396
rect 1344 42310 19838 42362
rect 19890 42310 19942 42362
rect 19994 42310 20046 42362
rect 20098 42310 50558 42362
rect 50610 42310 50662 42362
rect 50714 42310 50766 42362
rect 50818 42310 58576 42362
rect 1344 42276 58576 42310
rect 3502 42194 3554 42206
rect 16718 42194 16770 42206
rect 8866 42142 8878 42194
rect 8930 42142 8942 42194
rect 3502 42130 3554 42142
rect 16718 42130 16770 42142
rect 23662 42194 23714 42206
rect 23662 42130 23714 42142
rect 29374 42194 29426 42206
rect 35410 42142 35422 42194
rect 35474 42142 35486 42194
rect 29374 42130 29426 42142
rect 2270 42082 2322 42094
rect 2270 42018 2322 42030
rect 6414 42082 6466 42094
rect 17838 42082 17890 42094
rect 8978 42030 8990 42082
rect 9042 42030 9054 42082
rect 11106 42030 11118 42082
rect 11170 42030 11182 42082
rect 12114 42030 12126 42082
rect 12178 42030 12190 42082
rect 6414 42018 6466 42030
rect 17838 42018 17890 42030
rect 17950 42082 18002 42094
rect 30494 42082 30546 42094
rect 27906 42030 27918 42082
rect 27970 42030 27982 42082
rect 17950 42018 18002 42030
rect 30494 42018 30546 42030
rect 34526 42082 34578 42094
rect 34526 42018 34578 42030
rect 34974 42082 35026 42094
rect 41022 42082 41074 42094
rect 35186 42030 35198 42082
rect 35250 42030 35262 42082
rect 34974 42018 35026 42030
rect 41022 42018 41074 42030
rect 2494 41970 2546 41982
rect 2494 41906 2546 41918
rect 2718 41970 2770 41982
rect 2718 41906 2770 41918
rect 2830 41970 2882 41982
rect 2830 41906 2882 41918
rect 5294 41970 5346 41982
rect 16606 41970 16658 41982
rect 7410 41918 7422 41970
rect 7474 41918 7486 41970
rect 11442 41918 11454 41970
rect 11506 41918 11518 41970
rect 12226 41918 12238 41970
rect 12290 41918 12302 41970
rect 5294 41906 5346 41918
rect 16606 41906 16658 41918
rect 18174 41970 18226 41982
rect 18174 41906 18226 41918
rect 18622 41970 18674 41982
rect 18622 41906 18674 41918
rect 20190 41970 20242 41982
rect 20190 41906 20242 41918
rect 20414 41970 20466 41982
rect 20414 41906 20466 41918
rect 20638 41970 20690 41982
rect 20638 41906 20690 41918
rect 20862 41970 20914 41982
rect 20862 41906 20914 41918
rect 20974 41970 21026 41982
rect 20974 41906 21026 41918
rect 22094 41970 22146 41982
rect 22094 41906 22146 41918
rect 22206 41970 22258 41982
rect 22878 41970 22930 41982
rect 29934 41970 29986 41982
rect 22418 41918 22430 41970
rect 22482 41918 22494 41970
rect 29586 41918 29598 41970
rect 29650 41918 29662 41970
rect 22206 41906 22258 41918
rect 22878 41906 22930 41918
rect 29934 41906 29986 41918
rect 33518 41970 33570 41982
rect 35746 41918 35758 41970
rect 35810 41918 35822 41970
rect 33518 41906 33570 41918
rect 1822 41858 1874 41870
rect 1822 41794 1874 41806
rect 2606 41858 2658 41870
rect 2606 41794 2658 41806
rect 4062 41858 4114 41870
rect 19854 41858 19906 41870
rect 13010 41806 13022 41858
rect 13074 41806 13086 41858
rect 4062 41794 4114 41806
rect 19854 41794 19906 41806
rect 21534 41858 21586 41870
rect 21534 41794 21586 41806
rect 21870 41858 21922 41870
rect 21870 41794 21922 41806
rect 23214 41858 23266 41870
rect 23214 41794 23266 41806
rect 24670 41858 24722 41870
rect 24670 41794 24722 41806
rect 25342 41858 25394 41870
rect 25342 41794 25394 41806
rect 26574 41858 26626 41870
rect 26574 41794 26626 41806
rect 27246 41858 27298 41870
rect 27246 41794 27298 41806
rect 34078 41858 34130 41870
rect 34078 41794 34130 41806
rect 36206 41858 36258 41870
rect 36206 41794 36258 41806
rect 39902 41858 39954 41870
rect 39902 41794 39954 41806
rect 16718 41746 16770 41758
rect 16718 41682 16770 41694
rect 18510 41746 18562 41758
rect 18510 41682 18562 41694
rect 18846 41746 18898 41758
rect 18846 41682 18898 41694
rect 18958 41746 19010 41758
rect 18958 41682 19010 41694
rect 34302 41746 34354 41758
rect 34302 41682 34354 41694
rect 34638 41746 34690 41758
rect 34638 41682 34690 41694
rect 35422 41746 35474 41758
rect 35422 41682 35474 41694
rect 40910 41746 40962 41758
rect 40910 41682 40962 41694
rect 1344 41578 58576 41612
rect 1344 41526 4478 41578
rect 4530 41526 4582 41578
rect 4634 41526 4686 41578
rect 4738 41526 35198 41578
rect 35250 41526 35302 41578
rect 35354 41526 35406 41578
rect 35458 41526 58576 41578
rect 1344 41492 58576 41526
rect 13806 41410 13858 41422
rect 13806 41346 13858 41358
rect 14254 41410 14306 41422
rect 14254 41346 14306 41358
rect 21758 41410 21810 41422
rect 21758 41346 21810 41358
rect 22094 41410 22146 41422
rect 30046 41410 30098 41422
rect 28242 41358 28254 41410
rect 28306 41358 28318 41410
rect 35298 41358 35310 41410
rect 35362 41358 35374 41410
rect 22094 41346 22146 41358
rect 30046 41346 30098 41358
rect 7646 41298 7698 41310
rect 35982 41298 36034 41310
rect 9538 41246 9550 41298
rect 9602 41246 9614 41298
rect 12562 41246 12574 41298
rect 12626 41246 12638 41298
rect 18386 41246 18398 41298
rect 18450 41246 18462 41298
rect 24546 41246 24558 41298
rect 24610 41246 24622 41298
rect 27906 41246 27918 41298
rect 27970 41246 27982 41298
rect 7646 41234 7698 41246
rect 35982 41234 36034 41246
rect 1710 41186 1762 41198
rect 10334 41186 10386 41198
rect 5842 41134 5854 41186
rect 5906 41134 5918 41186
rect 9090 41134 9102 41186
rect 9154 41134 9166 41186
rect 9314 41134 9326 41186
rect 9378 41134 9390 41186
rect 1710 41122 1762 41134
rect 10334 41122 10386 41134
rect 10894 41186 10946 41198
rect 14030 41186 14082 41198
rect 19630 41186 19682 41198
rect 11890 41134 11902 41186
rect 11954 41134 11966 41186
rect 17154 41134 17166 41186
rect 17218 41134 17230 41186
rect 17602 41134 17614 41186
rect 17666 41134 17678 41186
rect 10894 41122 10946 41134
rect 14030 41122 14082 41134
rect 19630 41122 19682 41134
rect 19966 41186 20018 41198
rect 19966 41122 20018 41134
rect 20862 41186 20914 41198
rect 20862 41122 20914 41134
rect 21422 41186 21474 41198
rect 21422 41122 21474 41134
rect 21534 41186 21586 41198
rect 21534 41122 21586 41134
rect 21982 41186 22034 41198
rect 26910 41186 26962 41198
rect 29150 41186 29202 41198
rect 23314 41134 23326 41186
rect 23378 41134 23390 41186
rect 24882 41134 24894 41186
rect 24946 41134 24958 41186
rect 27122 41134 27134 41186
rect 27186 41134 27198 41186
rect 28354 41134 28366 41186
rect 28418 41134 28430 41186
rect 21982 41122 22034 41134
rect 26910 41122 26962 41134
rect 29150 41122 29202 41134
rect 29374 41186 29426 41198
rect 29374 41122 29426 41134
rect 29598 41186 29650 41198
rect 32958 41186 33010 41198
rect 34750 41186 34802 41198
rect 31266 41134 31278 41186
rect 31330 41134 31342 41186
rect 33506 41134 33518 41186
rect 33570 41134 33582 41186
rect 35298 41134 35310 41186
rect 35362 41134 35374 41186
rect 29598 41122 29650 41134
rect 32958 41122 33010 41134
rect 34750 41122 34802 41134
rect 2046 41074 2098 41086
rect 2046 41010 2098 41022
rect 2382 41074 2434 41086
rect 2382 41010 2434 41022
rect 2718 41074 2770 41086
rect 2718 41010 2770 41022
rect 6414 41074 6466 41086
rect 13582 41074 13634 41086
rect 18734 41074 18786 41086
rect 12114 41022 12126 41074
rect 12178 41022 12190 41074
rect 15698 41022 15710 41074
rect 15762 41022 15774 41074
rect 6414 41010 6466 41022
rect 13582 41010 13634 41022
rect 18734 41010 18786 41022
rect 19854 41074 19906 41086
rect 19854 41010 19906 41022
rect 20526 41074 20578 41086
rect 35870 41074 35922 41086
rect 23874 41022 23886 41074
rect 23938 41022 23950 41074
rect 25106 41022 25118 41074
rect 25170 41022 25182 41074
rect 31042 41022 31054 41074
rect 31106 41022 31118 41074
rect 34962 41022 34974 41074
rect 35026 41022 35038 41074
rect 20526 41010 20578 41022
rect 35870 41010 35922 41022
rect 14702 40962 14754 40974
rect 7858 40910 7870 40962
rect 7922 40910 7934 40962
rect 9538 40910 9550 40962
rect 9602 40910 9614 40962
rect 14702 40898 14754 40910
rect 15038 40962 15090 40974
rect 15038 40898 15090 40910
rect 20638 40962 20690 40974
rect 20638 40898 20690 40910
rect 22542 40962 22594 40974
rect 22542 40898 22594 40910
rect 22990 40962 23042 40974
rect 22990 40898 23042 40910
rect 30382 40962 30434 40974
rect 36094 40962 36146 40974
rect 33058 40910 33070 40962
rect 33122 40910 33134 40962
rect 35186 40910 35198 40962
rect 35250 40910 35262 40962
rect 30382 40898 30434 40910
rect 36094 40898 36146 40910
rect 1344 40794 58576 40828
rect 1344 40742 19838 40794
rect 19890 40742 19942 40794
rect 19994 40742 20046 40794
rect 20098 40742 50558 40794
rect 50610 40742 50662 40794
rect 50714 40742 50766 40794
rect 50818 40742 58576 40794
rect 1344 40708 58576 40742
rect 12238 40626 12290 40638
rect 12238 40562 12290 40574
rect 13022 40626 13074 40638
rect 18174 40626 18226 40638
rect 16370 40574 16382 40626
rect 16434 40574 16446 40626
rect 13022 40562 13074 40574
rect 18174 40562 18226 40574
rect 19518 40626 19570 40638
rect 19518 40562 19570 40574
rect 21086 40626 21138 40638
rect 21086 40562 21138 40574
rect 24110 40626 24162 40638
rect 27358 40626 27410 40638
rect 26674 40574 26686 40626
rect 26738 40574 26750 40626
rect 24110 40562 24162 40574
rect 27358 40562 27410 40574
rect 27694 40626 27746 40638
rect 27694 40562 27746 40574
rect 34078 40626 34130 40638
rect 34078 40562 34130 40574
rect 34526 40626 34578 40638
rect 34526 40562 34578 40574
rect 35758 40626 35810 40638
rect 35758 40562 35810 40574
rect 36318 40626 36370 40638
rect 36318 40562 36370 40574
rect 2046 40514 2098 40526
rect 2046 40450 2098 40462
rect 4174 40514 4226 40526
rect 4174 40450 4226 40462
rect 6190 40514 6242 40526
rect 11678 40514 11730 40526
rect 18734 40514 18786 40526
rect 9650 40462 9662 40514
rect 9714 40462 9726 40514
rect 15922 40462 15934 40514
rect 15986 40462 15998 40514
rect 16146 40462 16158 40514
rect 16210 40462 16222 40514
rect 17714 40462 17726 40514
rect 17778 40462 17790 40514
rect 6190 40450 6242 40462
rect 11678 40450 11730 40462
rect 18734 40450 18786 40462
rect 25230 40514 25282 40526
rect 25230 40450 25282 40462
rect 34974 40514 35026 40526
rect 37762 40462 37774 40514
rect 37826 40462 37838 40514
rect 34974 40450 35026 40462
rect 1710 40402 1762 40414
rect 1710 40338 1762 40350
rect 2494 40402 2546 40414
rect 2494 40338 2546 40350
rect 3390 40402 3442 40414
rect 5742 40402 5794 40414
rect 9102 40402 9154 40414
rect 11454 40402 11506 40414
rect 3602 40350 3614 40402
rect 3666 40350 3678 40402
rect 8082 40350 8094 40402
rect 8146 40350 8158 40402
rect 8418 40350 8430 40402
rect 8482 40350 8494 40402
rect 9874 40350 9886 40402
rect 9938 40350 9950 40402
rect 3390 40338 3442 40350
rect 5742 40338 5794 40350
rect 9102 40338 9154 40350
rect 11454 40338 11506 40350
rect 12798 40402 12850 40414
rect 15374 40402 15426 40414
rect 13346 40350 13358 40402
rect 13410 40350 13422 40402
rect 14354 40350 14366 40402
rect 14418 40350 14430 40402
rect 12798 40338 12850 40350
rect 15374 40338 15426 40350
rect 16606 40402 16658 40414
rect 18846 40402 18898 40414
rect 22542 40402 22594 40414
rect 35310 40402 35362 40414
rect 17490 40350 17502 40402
rect 17554 40350 17566 40402
rect 19058 40350 19070 40402
rect 19122 40350 19134 40402
rect 28578 40350 28590 40402
rect 28642 40350 28654 40402
rect 28802 40350 28814 40402
rect 28866 40350 28878 40402
rect 30146 40350 30158 40402
rect 30210 40350 30222 40402
rect 30818 40350 30830 40402
rect 30882 40350 30894 40402
rect 31378 40350 31390 40402
rect 31442 40350 31454 40402
rect 16606 40338 16658 40350
rect 18846 40338 18898 40350
rect 22542 40338 22594 40350
rect 35310 40338 35362 40350
rect 35422 40402 35474 40414
rect 35522 40350 35534 40402
rect 35586 40350 35598 40402
rect 36978 40350 36990 40402
rect 37042 40350 37054 40402
rect 35422 40338 35474 40350
rect 5406 40290 5458 40302
rect 11902 40290 11954 40302
rect 8754 40238 8766 40290
rect 8818 40238 8830 40290
rect 5406 40226 5458 40238
rect 11902 40226 11954 40238
rect 12910 40290 12962 40302
rect 12910 40226 12962 40238
rect 14814 40290 14866 40302
rect 14814 40226 14866 40238
rect 18510 40290 18562 40302
rect 18510 40226 18562 40238
rect 26126 40290 26178 40302
rect 30370 40238 30382 40290
rect 30434 40238 30446 40290
rect 34626 40238 34638 40290
rect 34690 40238 34702 40290
rect 39890 40238 39902 40290
rect 39954 40238 39966 40290
rect 26126 40226 26178 40238
rect 25342 40178 25394 40190
rect 25342 40114 25394 40126
rect 25566 40178 25618 40190
rect 25566 40114 25618 40126
rect 25678 40178 25730 40190
rect 25678 40114 25730 40126
rect 26350 40178 26402 40190
rect 26350 40114 26402 40126
rect 34302 40178 34354 40190
rect 34302 40114 34354 40126
rect 1344 40010 58576 40044
rect 1344 39958 4478 40010
rect 4530 39958 4582 40010
rect 4634 39958 4686 40010
rect 4738 39958 35198 40010
rect 35250 39958 35302 40010
rect 35354 39958 35406 40010
rect 35458 39958 58576 40010
rect 1344 39924 58576 39958
rect 27918 39842 27970 39854
rect 27918 39778 27970 39790
rect 28030 39842 28082 39854
rect 28030 39778 28082 39790
rect 28254 39842 28306 39854
rect 30258 39790 30270 39842
rect 30322 39790 30334 39842
rect 28254 39778 28306 39790
rect 20078 39730 20130 39742
rect 27582 39730 27634 39742
rect 8082 39678 8094 39730
rect 8146 39678 8158 39730
rect 11106 39678 11118 39730
rect 11170 39678 11182 39730
rect 22082 39678 22094 39730
rect 22146 39678 22158 39730
rect 26450 39678 26462 39730
rect 26514 39678 26526 39730
rect 20078 39666 20130 39678
rect 27582 39666 27634 39678
rect 29486 39730 29538 39742
rect 32162 39678 32174 39730
rect 32226 39678 32238 39730
rect 29486 39666 29538 39678
rect 16382 39618 16434 39630
rect 27022 39618 27074 39630
rect 30606 39618 30658 39630
rect 3938 39566 3950 39618
rect 4002 39566 4014 39618
rect 5058 39566 5070 39618
rect 5122 39566 5134 39618
rect 6738 39566 6750 39618
rect 6802 39566 6814 39618
rect 7970 39566 7982 39618
rect 8034 39566 8046 39618
rect 10546 39566 10558 39618
rect 10610 39566 10622 39618
rect 10770 39566 10782 39618
rect 10834 39566 10846 39618
rect 15026 39566 15038 39618
rect 15090 39566 15102 39618
rect 17378 39566 17390 39618
rect 17442 39566 17454 39618
rect 18946 39566 18958 39618
rect 19010 39566 19022 39618
rect 21298 39566 21310 39618
rect 21362 39566 21374 39618
rect 23314 39566 23326 39618
rect 23378 39566 23390 39618
rect 28466 39566 28478 39618
rect 28530 39566 28542 39618
rect 30034 39566 30046 39618
rect 30098 39566 30110 39618
rect 16382 39554 16434 39566
rect 27022 39554 27074 39566
rect 30606 39554 30658 39566
rect 30830 39618 30882 39630
rect 31490 39566 31502 39618
rect 31554 39566 31566 39618
rect 31714 39566 31726 39618
rect 31778 39566 31790 39618
rect 33954 39566 33966 39618
rect 34018 39566 34030 39618
rect 34290 39566 34302 39618
rect 34354 39566 34366 39618
rect 30830 39554 30882 39566
rect 2830 39506 2882 39518
rect 2830 39442 2882 39454
rect 3054 39506 3106 39518
rect 14702 39506 14754 39518
rect 23886 39506 23938 39518
rect 3378 39454 3390 39506
rect 3442 39454 3454 39506
rect 4946 39454 4958 39506
rect 5010 39454 5022 39506
rect 7186 39454 7198 39506
rect 7250 39454 7262 39506
rect 8194 39454 8206 39506
rect 8258 39454 8270 39506
rect 18162 39454 18174 39506
rect 18226 39454 18238 39506
rect 27122 39454 27134 39506
rect 27186 39454 27198 39506
rect 33730 39454 33742 39506
rect 33794 39454 33806 39506
rect 34626 39454 34638 39506
rect 34690 39454 34702 39506
rect 3054 39442 3106 39454
rect 14702 39442 14754 39454
rect 23886 39442 23938 39454
rect 2942 39394 2994 39406
rect 6078 39394 6130 39406
rect 14142 39394 14194 39406
rect 19518 39394 19570 39406
rect 3490 39342 3502 39394
rect 3554 39342 3566 39394
rect 10994 39342 11006 39394
rect 11058 39342 11070 39394
rect 15138 39342 15150 39394
rect 15202 39342 15214 39394
rect 2942 39330 2994 39342
rect 6078 39330 6130 39342
rect 14142 39330 14194 39342
rect 19518 39330 19570 39342
rect 22990 39394 23042 39406
rect 22990 39330 23042 39342
rect 1344 39226 58576 39260
rect 1344 39174 19838 39226
rect 19890 39174 19942 39226
rect 19994 39174 20046 39226
rect 20098 39174 50558 39226
rect 50610 39174 50662 39226
rect 50714 39174 50766 39226
rect 50818 39174 58576 39226
rect 1344 39140 58576 39174
rect 5294 39058 5346 39070
rect 11790 39058 11842 39070
rect 15038 39058 15090 39070
rect 5842 39006 5854 39058
rect 5906 39006 5918 39058
rect 13010 39006 13022 39058
rect 13074 39006 13086 39058
rect 5294 38994 5346 39006
rect 11790 38994 11842 39006
rect 15038 38994 15090 39006
rect 15262 39058 15314 39070
rect 15262 38994 15314 39006
rect 19406 39058 19458 39070
rect 19406 38994 19458 39006
rect 22206 39058 22258 39070
rect 22206 38994 22258 39006
rect 25118 39058 25170 39070
rect 25118 38994 25170 39006
rect 27582 39058 27634 39070
rect 27582 38994 27634 39006
rect 28702 39058 28754 39070
rect 28702 38994 28754 39006
rect 29262 39058 29314 39070
rect 29262 38994 29314 39006
rect 21310 38946 21362 38958
rect 2370 38894 2382 38946
rect 2434 38894 2446 38946
rect 3490 38894 3502 38946
rect 3554 38894 3566 38946
rect 5730 38894 5742 38946
rect 5794 38894 5806 38946
rect 7298 38894 7310 38946
rect 7362 38894 7374 38946
rect 21310 38882 21362 38894
rect 24222 38946 24274 38958
rect 27918 38946 27970 38958
rect 26674 38894 26686 38946
rect 26738 38894 26750 38946
rect 24222 38882 24274 38894
rect 27918 38882 27970 38894
rect 30942 38946 30994 38958
rect 32386 38894 32398 38946
rect 32450 38894 32462 38946
rect 34402 38894 34414 38946
rect 34466 38894 34478 38946
rect 35298 38894 35310 38946
rect 35362 38894 35374 38946
rect 38210 38894 38222 38946
rect 38274 38894 38286 38946
rect 30942 38882 30994 38894
rect 3838 38834 3890 38846
rect 2594 38782 2606 38834
rect 2658 38782 2670 38834
rect 3838 38770 3890 38782
rect 4286 38834 4338 38846
rect 6750 38834 6802 38846
rect 5618 38782 5630 38834
rect 5682 38782 5694 38834
rect 4286 38770 4338 38782
rect 6750 38770 6802 38782
rect 7758 38834 7810 38846
rect 7758 38770 7810 38782
rect 7982 38834 8034 38846
rect 7982 38770 8034 38782
rect 12350 38834 12402 38846
rect 13918 38834 13970 38846
rect 12786 38782 12798 38834
rect 12850 38782 12862 38834
rect 12350 38770 12402 38782
rect 13918 38770 13970 38782
rect 14478 38834 14530 38846
rect 14478 38770 14530 38782
rect 14814 38834 14866 38846
rect 14814 38770 14866 38782
rect 15486 38834 15538 38846
rect 15486 38770 15538 38782
rect 21198 38834 21250 38846
rect 21982 38834 22034 38846
rect 21522 38782 21534 38834
rect 21586 38782 21598 38834
rect 21198 38770 21250 38782
rect 21982 38770 22034 38782
rect 23774 38834 23826 38846
rect 23774 38770 23826 38782
rect 24670 38834 24722 38846
rect 24670 38770 24722 38782
rect 25790 38834 25842 38846
rect 25790 38770 25842 38782
rect 26014 38834 26066 38846
rect 26014 38770 26066 38782
rect 26910 38834 26962 38846
rect 27122 38782 27134 38834
rect 27186 38782 27198 38834
rect 31154 38782 31166 38834
rect 31218 38782 31230 38834
rect 31714 38782 31726 38834
rect 31778 38782 31790 38834
rect 32498 38782 32510 38834
rect 32562 38782 32574 38834
rect 34290 38782 34302 38834
rect 34354 38782 34366 38834
rect 36754 38782 36766 38834
rect 36818 38782 36830 38834
rect 37426 38782 37438 38834
rect 37490 38782 37502 38834
rect 26910 38770 26962 38782
rect 1822 38722 1874 38734
rect 1822 38658 1874 38670
rect 8094 38722 8146 38734
rect 8094 38658 8146 38670
rect 8654 38722 8706 38734
rect 8654 38658 8706 38670
rect 16270 38722 16322 38734
rect 16270 38658 16322 38670
rect 18062 38722 18114 38734
rect 18062 38658 18114 38670
rect 18622 38722 18674 38734
rect 18622 38658 18674 38670
rect 19070 38722 19122 38734
rect 19070 38658 19122 38670
rect 20302 38722 20354 38734
rect 20302 38658 20354 38670
rect 20974 38722 21026 38734
rect 20974 38658 21026 38670
rect 22766 38722 22818 38734
rect 22766 38658 22818 38670
rect 23214 38722 23266 38734
rect 25566 38722 25618 38734
rect 24546 38719 24558 38722
rect 23214 38658 23266 38670
rect 24337 38673 24558 38719
rect 7646 38610 7698 38622
rect 7646 38546 7698 38558
rect 15374 38610 15426 38622
rect 23986 38558 23998 38610
rect 24050 38607 24062 38610
rect 24337 38607 24383 38673
rect 24546 38670 24558 38673
rect 24610 38670 24622 38722
rect 25566 38658 25618 38670
rect 26238 38722 26290 38734
rect 26238 38658 26290 38670
rect 26574 38722 26626 38734
rect 33618 38670 33630 38722
rect 33682 38670 33694 38722
rect 40338 38670 40350 38722
rect 40402 38670 40414 38722
rect 26574 38658 26626 38670
rect 24050 38561 24383 38607
rect 24050 38558 24062 38561
rect 15374 38546 15426 38558
rect 1344 38442 58576 38476
rect 1344 38390 4478 38442
rect 4530 38390 4582 38442
rect 4634 38390 4686 38442
rect 4738 38390 35198 38442
rect 35250 38390 35302 38442
rect 35354 38390 35406 38442
rect 35458 38390 58576 38442
rect 1344 38356 58576 38390
rect 4958 38274 5010 38286
rect 4958 38210 5010 38222
rect 11230 38274 11282 38286
rect 19070 38274 19122 38286
rect 16594 38271 16606 38274
rect 11230 38210 11282 38222
rect 16161 38225 16606 38271
rect 3950 38162 4002 38174
rect 13358 38162 13410 38174
rect 7410 38110 7422 38162
rect 7474 38110 7486 38162
rect 12226 38110 12238 38162
rect 12290 38110 12302 38162
rect 15138 38110 15150 38162
rect 15202 38110 15214 38162
rect 3950 38098 4002 38110
rect 13358 38098 13410 38110
rect 2494 38050 2546 38062
rect 2494 37986 2546 37998
rect 3054 38050 3106 38062
rect 3054 37986 3106 37998
rect 3614 38050 3666 38062
rect 3614 37986 3666 37998
rect 4734 38050 4786 38062
rect 4734 37986 4786 37998
rect 5630 38050 5682 38062
rect 9214 38050 9266 38062
rect 6514 37998 6526 38050
rect 6578 37998 6590 38050
rect 7522 37998 7534 38050
rect 7586 37998 7598 38050
rect 5630 37986 5682 37998
rect 9214 37986 9266 37998
rect 9550 38050 9602 38062
rect 11790 38050 11842 38062
rect 9986 37998 9998 38050
rect 10050 37998 10062 38050
rect 9550 37986 9602 37998
rect 11790 37986 11842 37998
rect 11902 38050 11954 38062
rect 14030 38050 14082 38062
rect 12338 37998 12350 38050
rect 12402 37998 12414 38050
rect 15026 37998 15038 38050
rect 15090 37998 15102 38050
rect 15586 37998 15598 38050
rect 15650 37998 15662 38050
rect 11902 37986 11954 37998
rect 14030 37986 14082 37998
rect 1710 37938 1762 37950
rect 1710 37874 1762 37886
rect 2606 37938 2658 37950
rect 4286 37938 4338 37950
rect 10894 37938 10946 37950
rect 4050 37886 4062 37938
rect 4114 37886 4126 37938
rect 6738 37886 6750 37938
rect 6802 37886 6814 37938
rect 2606 37874 2658 37886
rect 4286 37874 4338 37886
rect 10894 37874 10946 37886
rect 11342 37938 11394 37950
rect 11342 37874 11394 37886
rect 13470 37938 13522 37950
rect 14466 37886 14478 37938
rect 14530 37886 14542 37938
rect 15922 37886 15934 37938
rect 15986 37935 15998 37938
rect 16161 37935 16207 38225
rect 16594 38222 16606 38225
rect 16658 38222 16670 38274
rect 19070 38210 19122 38222
rect 20638 38274 20690 38286
rect 20638 38210 20690 38222
rect 37774 38274 37826 38286
rect 37774 38210 37826 38222
rect 19630 38162 19682 38174
rect 19630 38098 19682 38110
rect 22878 38162 22930 38174
rect 28366 38162 28418 38174
rect 26226 38110 26238 38162
rect 26290 38110 26302 38162
rect 22878 38098 22930 38110
rect 28366 38098 28418 38110
rect 30046 38162 30098 38174
rect 30046 38098 30098 38110
rect 32846 38162 32898 38174
rect 36430 38162 36482 38174
rect 34178 38110 34190 38162
rect 34242 38110 34254 38162
rect 37202 38110 37214 38162
rect 37266 38110 37278 38162
rect 32846 38098 32898 38110
rect 36430 38098 36482 38110
rect 17166 38050 17218 38062
rect 17166 37986 17218 37998
rect 17838 38050 17890 38062
rect 18510 38050 18562 38062
rect 18274 37998 18286 38050
rect 18338 37998 18350 38050
rect 17838 37986 17890 37998
rect 18510 37986 18562 37998
rect 18734 38050 18786 38062
rect 18734 37986 18786 37998
rect 18958 38050 19010 38062
rect 18958 37986 19010 37998
rect 19966 38050 20018 38062
rect 29822 38050 29874 38062
rect 20290 37998 20302 38050
rect 20354 37998 20366 38050
rect 24098 37998 24110 38050
rect 24162 37998 24174 38050
rect 26114 37998 26126 38050
rect 26178 37998 26190 38050
rect 28578 37998 28590 38050
rect 28642 37998 28654 38050
rect 19966 37986 20018 37998
rect 29822 37986 29874 37998
rect 30494 38050 30546 38062
rect 30494 37986 30546 37998
rect 31838 38050 31890 38062
rect 37998 38050 38050 38062
rect 33282 37998 33294 38050
rect 33346 37998 33358 38050
rect 31838 37986 31890 37998
rect 37998 37986 38050 37998
rect 38222 38050 38274 38062
rect 38222 37986 38274 37998
rect 38446 38050 38498 38062
rect 38446 37986 38498 37998
rect 15986 37889 16207 37935
rect 17726 37938 17778 37950
rect 27246 37938 27298 37950
rect 15986 37886 15998 37889
rect 19730 37886 19742 37938
rect 19794 37886 19806 37938
rect 24210 37886 24222 37938
rect 24274 37886 24286 37938
rect 13470 37874 13522 37886
rect 17726 37874 17778 37886
rect 27246 37874 27298 37886
rect 28254 37938 28306 37950
rect 28254 37874 28306 37886
rect 30606 37938 30658 37950
rect 30606 37874 30658 37886
rect 32062 37938 32114 37950
rect 32062 37874 32114 37886
rect 32174 37938 32226 37950
rect 32174 37874 32226 37886
rect 2046 37826 2098 37838
rect 2046 37762 2098 37774
rect 2830 37826 2882 37838
rect 2830 37762 2882 37774
rect 6190 37826 6242 37838
rect 10670 37826 10722 37838
rect 6850 37774 6862 37826
rect 6914 37774 6926 37826
rect 6190 37762 6242 37774
rect 10670 37762 10722 37774
rect 11118 37826 11170 37838
rect 11118 37762 11170 37774
rect 12126 37826 12178 37838
rect 12126 37762 12178 37774
rect 12798 37826 12850 37838
rect 12798 37762 12850 37774
rect 13694 37826 13746 37838
rect 13694 37762 13746 37774
rect 13918 37826 13970 37838
rect 13918 37762 13970 37774
rect 15710 37826 15762 37838
rect 15710 37762 15762 37774
rect 16382 37826 16434 37838
rect 16382 37762 16434 37774
rect 17278 37826 17330 37838
rect 17278 37762 17330 37774
rect 17502 37826 17554 37838
rect 17502 37762 17554 37774
rect 21534 37826 21586 37838
rect 21534 37762 21586 37774
rect 21982 37826 22034 37838
rect 21982 37762 22034 37774
rect 22542 37826 22594 37838
rect 22542 37762 22594 37774
rect 23438 37826 23490 37838
rect 23438 37762 23490 37774
rect 23774 37826 23826 37838
rect 23774 37762 23826 37774
rect 29710 37826 29762 37838
rect 29710 37762 29762 37774
rect 33742 37826 33794 37838
rect 33742 37762 33794 37774
rect 1344 37658 58576 37692
rect 1344 37606 19838 37658
rect 19890 37606 19942 37658
rect 19994 37606 20046 37658
rect 20098 37606 50558 37658
rect 50610 37606 50662 37658
rect 50714 37606 50766 37658
rect 50818 37606 58576 37658
rect 1344 37572 58576 37606
rect 2606 37490 2658 37502
rect 2606 37426 2658 37438
rect 2830 37490 2882 37502
rect 2830 37426 2882 37438
rect 6302 37490 6354 37502
rect 10558 37490 10610 37502
rect 8194 37438 8206 37490
rect 8258 37438 8270 37490
rect 6302 37426 6354 37438
rect 10558 37426 10610 37438
rect 12574 37490 12626 37502
rect 12574 37426 12626 37438
rect 13022 37490 13074 37502
rect 13022 37426 13074 37438
rect 18622 37490 18674 37502
rect 18622 37426 18674 37438
rect 19182 37490 19234 37502
rect 19182 37426 19234 37438
rect 19406 37490 19458 37502
rect 19406 37426 19458 37438
rect 25230 37490 25282 37502
rect 26798 37490 26850 37502
rect 26002 37438 26014 37490
rect 26066 37438 26078 37490
rect 25230 37426 25282 37438
rect 26798 37426 26850 37438
rect 29598 37490 29650 37502
rect 29598 37426 29650 37438
rect 29710 37490 29762 37502
rect 29710 37426 29762 37438
rect 32062 37490 32114 37502
rect 32062 37426 32114 37438
rect 39902 37490 39954 37502
rect 39902 37426 39954 37438
rect 2046 37378 2098 37390
rect 2046 37314 2098 37326
rect 2494 37378 2546 37390
rect 2494 37314 2546 37326
rect 9774 37378 9826 37390
rect 15822 37378 15874 37390
rect 12114 37326 12126 37378
rect 12178 37326 12190 37378
rect 9774 37314 9826 37326
rect 15822 37314 15874 37326
rect 16494 37378 16546 37390
rect 18286 37378 18338 37390
rect 17826 37326 17838 37378
rect 17890 37326 17902 37378
rect 16494 37314 16546 37326
rect 18286 37314 18338 37326
rect 18398 37378 18450 37390
rect 25454 37378 25506 37390
rect 21186 37326 21198 37378
rect 21250 37326 21262 37378
rect 18398 37314 18450 37326
rect 25454 37314 25506 37326
rect 25566 37378 25618 37390
rect 29038 37378 29090 37390
rect 26226 37326 26238 37378
rect 26290 37326 26302 37378
rect 25566 37314 25618 37326
rect 29038 37314 29090 37326
rect 29486 37378 29538 37390
rect 40238 37378 40290 37390
rect 35858 37326 35870 37378
rect 35922 37326 35934 37378
rect 39554 37326 39566 37378
rect 39618 37326 39630 37378
rect 29486 37314 29538 37326
rect 40238 37314 40290 37326
rect 1710 37266 1762 37278
rect 8654 37266 8706 37278
rect 7746 37214 7758 37266
rect 7810 37214 7822 37266
rect 1710 37202 1762 37214
rect 8654 37202 8706 37214
rect 8766 37266 8818 37278
rect 9662 37266 9714 37278
rect 8978 37214 8990 37266
rect 9042 37214 9054 37266
rect 8766 37202 8818 37214
rect 9662 37202 9714 37214
rect 9886 37266 9938 37278
rect 15150 37266 15202 37278
rect 10098 37214 10110 37266
rect 10162 37214 10174 37266
rect 11890 37214 11902 37266
rect 11954 37214 11966 37266
rect 9886 37202 9938 37214
rect 15150 37202 15202 37214
rect 15374 37266 15426 37278
rect 17502 37266 17554 37278
rect 16034 37214 16046 37266
rect 16098 37214 16110 37266
rect 16258 37214 16270 37266
rect 16322 37214 16334 37266
rect 15374 37202 15426 37214
rect 17502 37202 17554 37214
rect 19070 37266 19122 37278
rect 27694 37266 27746 37278
rect 20066 37214 20078 37266
rect 20130 37214 20142 37266
rect 22642 37214 22654 37266
rect 22706 37214 22718 37266
rect 22866 37214 22878 37266
rect 22930 37214 22942 37266
rect 23202 37214 23214 37266
rect 23266 37214 23278 37266
rect 23538 37214 23550 37266
rect 23602 37214 23614 37266
rect 26562 37214 26574 37266
rect 26626 37214 26638 37266
rect 19070 37202 19122 37214
rect 27694 37202 27746 37214
rect 29822 37266 29874 37278
rect 32286 37266 32338 37278
rect 30034 37214 30046 37266
rect 30098 37214 30110 37266
rect 31042 37214 31054 37266
rect 31106 37214 31118 37266
rect 31266 37214 31278 37266
rect 31330 37214 31342 37266
rect 31490 37214 31502 37266
rect 31554 37214 31566 37266
rect 29822 37202 29874 37214
rect 32286 37202 32338 37214
rect 34190 37266 34242 37278
rect 34190 37202 34242 37214
rect 34750 37266 34802 37278
rect 35074 37214 35086 37266
rect 35138 37214 35150 37266
rect 38658 37214 38670 37266
rect 38722 37214 38734 37266
rect 34750 37202 34802 37214
rect 3166 37154 3218 37166
rect 14926 37154 14978 37166
rect 7410 37102 7422 37154
rect 7474 37102 7486 37154
rect 3166 37090 3218 37102
rect 14926 37090 14978 37102
rect 16158 37154 16210 37166
rect 16158 37090 16210 37102
rect 21422 37154 21474 37166
rect 21422 37090 21474 37102
rect 27246 37154 27298 37166
rect 27246 37090 27298 37102
rect 27918 37154 27970 37166
rect 27918 37090 27970 37102
rect 28478 37154 28530 37166
rect 37998 37154 38050 37166
rect 31938 37102 31950 37154
rect 32002 37102 32014 37154
rect 28478 37090 28530 37102
rect 37998 37090 38050 37102
rect 39118 37154 39170 37166
rect 39118 37090 39170 37102
rect 27470 37042 27522 37054
rect 40350 37042 40402 37054
rect 30482 36990 30494 37042
rect 30546 36990 30558 37042
rect 27470 36978 27522 36990
rect 40350 36978 40402 36990
rect 1344 36874 58576 36908
rect 1344 36822 4478 36874
rect 4530 36822 4582 36874
rect 4634 36822 4686 36874
rect 4738 36822 35198 36874
rect 35250 36822 35302 36874
rect 35354 36822 35406 36874
rect 35458 36822 58576 36874
rect 1344 36788 58576 36822
rect 14142 36706 14194 36718
rect 14142 36642 14194 36654
rect 7982 36594 8034 36606
rect 3602 36542 3614 36594
rect 3666 36542 3678 36594
rect 7074 36542 7086 36594
rect 7138 36542 7150 36594
rect 7982 36530 8034 36542
rect 8206 36594 8258 36606
rect 8206 36530 8258 36542
rect 12910 36594 12962 36606
rect 19294 36594 19346 36606
rect 18050 36542 18062 36594
rect 18114 36542 18126 36594
rect 12910 36530 12962 36542
rect 19294 36530 19346 36542
rect 19854 36594 19906 36606
rect 19854 36530 19906 36542
rect 27582 36594 27634 36606
rect 27582 36530 27634 36542
rect 31726 36594 31778 36606
rect 37314 36542 37326 36594
rect 37378 36542 37390 36594
rect 39330 36542 39342 36594
rect 39394 36542 39406 36594
rect 31726 36530 31778 36542
rect 8654 36482 8706 36494
rect 2482 36430 2494 36482
rect 2546 36430 2558 36482
rect 2706 36430 2718 36482
rect 2770 36430 2782 36482
rect 3266 36430 3278 36482
rect 3330 36430 3342 36482
rect 5730 36430 5742 36482
rect 5794 36430 5806 36482
rect 8654 36418 8706 36430
rect 14366 36482 14418 36494
rect 14366 36418 14418 36430
rect 20414 36482 20466 36494
rect 20414 36418 20466 36430
rect 20750 36482 20802 36494
rect 28702 36482 28754 36494
rect 22530 36430 22542 36482
rect 22594 36430 22606 36482
rect 24210 36430 24222 36482
rect 24274 36430 24286 36482
rect 25330 36430 25342 36482
rect 25394 36430 25406 36482
rect 25778 36430 25790 36482
rect 25842 36430 25854 36482
rect 26002 36430 26014 36482
rect 26066 36430 26078 36482
rect 20750 36418 20802 36430
rect 28702 36418 28754 36430
rect 32734 36482 32786 36494
rect 34414 36482 34466 36494
rect 33170 36430 33182 36482
rect 33234 36430 33246 36482
rect 36194 36430 36206 36482
rect 36258 36430 36270 36482
rect 37986 36430 37998 36482
rect 38050 36430 38062 36482
rect 38546 36430 38558 36482
rect 38610 36430 38622 36482
rect 32734 36418 32786 36430
rect 34414 36418 34466 36430
rect 6750 36370 6802 36382
rect 1922 36318 1934 36370
rect 1986 36318 1998 36370
rect 3826 36318 3838 36370
rect 3890 36318 3902 36370
rect 5954 36318 5966 36370
rect 6018 36318 6030 36370
rect 6750 36306 6802 36318
rect 13806 36370 13858 36382
rect 13806 36306 13858 36318
rect 17502 36370 17554 36382
rect 17502 36306 17554 36318
rect 18062 36370 18114 36382
rect 18062 36306 18114 36318
rect 18286 36370 18338 36382
rect 28366 36370 28418 36382
rect 22978 36318 22990 36370
rect 23042 36318 23054 36370
rect 18286 36306 18338 36318
rect 28366 36306 28418 36318
rect 35646 36370 35698 36382
rect 35646 36306 35698 36318
rect 4286 36258 4338 36270
rect 4286 36194 4338 36206
rect 4846 36258 4898 36270
rect 4846 36194 4898 36206
rect 8990 36258 9042 36270
rect 8990 36194 9042 36206
rect 10558 36258 10610 36270
rect 10558 36194 10610 36206
rect 14030 36258 14082 36270
rect 14030 36194 14082 36206
rect 17838 36258 17890 36270
rect 17838 36194 17890 36206
rect 18958 36258 19010 36270
rect 18958 36194 19010 36206
rect 20302 36258 20354 36270
rect 20302 36194 20354 36206
rect 20638 36258 20690 36270
rect 20638 36194 20690 36206
rect 21534 36258 21586 36270
rect 21534 36194 21586 36206
rect 21870 36258 21922 36270
rect 28030 36258 28082 36270
rect 23874 36206 23886 36258
rect 23938 36206 23950 36258
rect 21870 36194 21922 36206
rect 28030 36194 28082 36206
rect 28478 36258 28530 36270
rect 28478 36194 28530 36206
rect 29262 36258 29314 36270
rect 29262 36194 29314 36206
rect 29710 36258 29762 36270
rect 29710 36194 29762 36206
rect 32286 36258 32338 36270
rect 32286 36194 32338 36206
rect 33854 36258 33906 36270
rect 33854 36194 33906 36206
rect 40126 36258 40178 36270
rect 40126 36194 40178 36206
rect 40910 36258 40962 36270
rect 40910 36194 40962 36206
rect 1344 36090 58576 36124
rect 1344 36038 19838 36090
rect 19890 36038 19942 36090
rect 19994 36038 20046 36090
rect 20098 36038 50558 36090
rect 50610 36038 50662 36090
rect 50714 36038 50766 36090
rect 50818 36038 58576 36090
rect 1344 36004 58576 36038
rect 2494 35922 2546 35934
rect 2494 35858 2546 35870
rect 3502 35922 3554 35934
rect 3502 35858 3554 35870
rect 4622 35922 4674 35934
rect 4622 35858 4674 35870
rect 5742 35922 5794 35934
rect 5742 35858 5794 35870
rect 7646 35922 7698 35934
rect 7646 35858 7698 35870
rect 10110 35922 10162 35934
rect 10110 35858 10162 35870
rect 10446 35922 10498 35934
rect 10446 35858 10498 35870
rect 12014 35922 12066 35934
rect 12014 35858 12066 35870
rect 12574 35922 12626 35934
rect 12574 35858 12626 35870
rect 15038 35922 15090 35934
rect 19742 35922 19794 35934
rect 28254 35922 28306 35934
rect 19058 35870 19070 35922
rect 19122 35870 19134 35922
rect 20850 35870 20862 35922
rect 20914 35870 20926 35922
rect 27458 35870 27470 35922
rect 27522 35870 27534 35922
rect 15038 35858 15090 35870
rect 19742 35858 19794 35870
rect 28254 35858 28306 35870
rect 28478 35922 28530 35934
rect 40350 35922 40402 35934
rect 33394 35870 33406 35922
rect 33458 35870 33470 35922
rect 28478 35858 28530 35870
rect 40350 35858 40402 35870
rect 40910 35922 40962 35934
rect 40910 35858 40962 35870
rect 2270 35810 2322 35822
rect 2270 35746 2322 35758
rect 3726 35810 3778 35822
rect 3726 35746 3778 35758
rect 10334 35810 10386 35822
rect 10334 35746 10386 35758
rect 14814 35810 14866 35822
rect 19966 35810 20018 35822
rect 33854 35810 33906 35822
rect 17714 35758 17726 35810
rect 17778 35758 17790 35810
rect 19282 35758 19294 35810
rect 19346 35758 19358 35810
rect 20514 35758 20526 35810
rect 20578 35758 20590 35810
rect 22866 35758 22878 35810
rect 22930 35758 22942 35810
rect 23874 35758 23886 35810
rect 23938 35758 23950 35810
rect 25442 35758 25454 35810
rect 25506 35758 25518 35810
rect 14814 35746 14866 35758
rect 19966 35746 20018 35758
rect 33854 35746 33906 35758
rect 36430 35810 36482 35822
rect 39230 35810 39282 35822
rect 37426 35758 37438 35810
rect 37490 35758 37502 35810
rect 37650 35758 37662 35810
rect 37714 35758 37726 35810
rect 36430 35746 36482 35758
rect 39230 35746 39282 35758
rect 2606 35698 2658 35710
rect 2606 35634 2658 35646
rect 2718 35698 2770 35710
rect 2718 35634 2770 35646
rect 2830 35698 2882 35710
rect 2830 35634 2882 35646
rect 3166 35698 3218 35710
rect 3166 35634 3218 35646
rect 9774 35698 9826 35710
rect 9774 35634 9826 35646
rect 12126 35698 12178 35710
rect 14702 35698 14754 35710
rect 18734 35698 18786 35710
rect 13906 35646 13918 35698
rect 13970 35646 13982 35698
rect 17602 35646 17614 35698
rect 17666 35646 17678 35698
rect 12126 35634 12178 35646
rect 14702 35634 14754 35646
rect 18734 35634 18786 35646
rect 20078 35698 20130 35710
rect 27806 35698 27858 35710
rect 20962 35646 20974 35698
rect 21026 35646 21038 35698
rect 22978 35646 22990 35698
rect 23042 35646 23054 35698
rect 23538 35646 23550 35698
rect 23602 35646 23614 35698
rect 25218 35646 25230 35698
rect 25282 35646 25294 35698
rect 20078 35634 20130 35646
rect 27806 35634 27858 35646
rect 28142 35698 28194 35710
rect 28142 35634 28194 35646
rect 28814 35698 28866 35710
rect 28814 35634 28866 35646
rect 34974 35698 35026 35710
rect 37090 35646 37102 35698
rect 37154 35646 37166 35698
rect 38546 35646 38558 35698
rect 38610 35646 38622 35698
rect 39666 35646 39678 35698
rect 39730 35646 39742 35698
rect 34974 35634 35026 35646
rect 6302 35586 6354 35598
rect 3490 35534 3502 35586
rect 3554 35534 3566 35586
rect 6302 35522 6354 35534
rect 8206 35586 8258 35598
rect 8206 35522 8258 35534
rect 10782 35586 10834 35598
rect 10782 35522 10834 35534
rect 11566 35586 11618 35598
rect 11566 35522 11618 35534
rect 13022 35586 13074 35598
rect 13022 35522 13074 35534
rect 14366 35586 14418 35598
rect 14366 35522 14418 35534
rect 15374 35586 15426 35598
rect 26686 35586 26738 35598
rect 23426 35534 23438 35586
rect 23490 35534 23502 35586
rect 25330 35534 25342 35586
rect 25394 35534 25406 35586
rect 15374 35522 15426 35534
rect 26686 35522 26738 35534
rect 27134 35586 27186 35598
rect 27134 35522 27186 35534
rect 29262 35586 29314 35598
rect 41346 35534 41358 35586
rect 41410 35534 41422 35586
rect 29262 35522 29314 35534
rect 12014 35474 12066 35486
rect 12014 35410 12066 35422
rect 1344 35306 58576 35340
rect 1344 35254 4478 35306
rect 4530 35254 4582 35306
rect 4634 35254 4686 35306
rect 4738 35254 35198 35306
rect 35250 35254 35302 35306
rect 35354 35254 35406 35306
rect 35458 35254 58576 35306
rect 1344 35220 58576 35254
rect 12350 35138 12402 35150
rect 12350 35074 12402 35086
rect 9886 35026 9938 35038
rect 18734 35026 18786 35038
rect 2818 34974 2830 35026
rect 2882 34974 2894 35026
rect 17266 34974 17278 35026
rect 17330 34974 17342 35026
rect 9886 34962 9938 34974
rect 18734 34962 18786 34974
rect 20302 35026 20354 35038
rect 20302 34962 20354 34974
rect 26462 35026 26514 35038
rect 26462 34962 26514 34974
rect 26798 35026 26850 35038
rect 26798 34962 26850 34974
rect 27694 35026 27746 35038
rect 29362 34974 29374 35026
rect 29426 34974 29438 35026
rect 30482 34974 30494 35026
rect 30546 34974 30558 35026
rect 27694 34962 27746 34974
rect 8094 34914 8146 34926
rect 6514 34862 6526 34914
rect 6578 34862 6590 34914
rect 8094 34850 8146 34862
rect 8654 34914 8706 34926
rect 8654 34850 8706 34862
rect 10446 34914 10498 34926
rect 10446 34850 10498 34862
rect 10894 34914 10946 34926
rect 12574 34914 12626 34926
rect 19406 34914 19458 34926
rect 12226 34862 12238 34914
rect 12290 34862 12302 34914
rect 13458 34862 13470 34914
rect 13522 34862 13534 34914
rect 14914 34862 14926 34914
rect 14978 34862 14990 34914
rect 16034 34862 16046 34914
rect 16098 34862 16110 34914
rect 16930 34862 16942 34914
rect 16994 34862 17006 34914
rect 10894 34850 10946 34862
rect 12574 34850 12626 34862
rect 19406 34850 19458 34862
rect 20862 34914 20914 34926
rect 26686 34914 26738 34926
rect 22866 34862 22878 34914
rect 22930 34862 22942 34914
rect 23762 34862 23774 34914
rect 23826 34862 23838 34914
rect 25218 34862 25230 34914
rect 25282 34862 25294 34914
rect 20862 34850 20914 34862
rect 26686 34850 26738 34862
rect 27022 34914 27074 34926
rect 27022 34850 27074 34862
rect 27134 34914 27186 34926
rect 27134 34850 27186 34862
rect 27582 34914 27634 34926
rect 27582 34850 27634 34862
rect 27806 34914 27858 34926
rect 27806 34850 27858 34862
rect 29822 34914 29874 34926
rect 29822 34850 29874 34862
rect 30942 34914 30994 34926
rect 30942 34850 30994 34862
rect 32398 34914 32450 34926
rect 32398 34850 32450 34862
rect 32734 34914 32786 34926
rect 35410 34862 35422 34914
rect 35474 34862 35486 34914
rect 36418 34862 36430 34914
rect 36482 34862 36494 34914
rect 38546 34862 38558 34914
rect 38610 34862 38622 34914
rect 38994 34862 39006 34914
rect 39058 34862 39070 34914
rect 32734 34850 32786 34862
rect 2270 34802 2322 34814
rect 2270 34738 2322 34750
rect 2718 34802 2770 34814
rect 2718 34738 2770 34750
rect 2830 34802 2882 34814
rect 2830 34738 2882 34750
rect 5630 34802 5682 34814
rect 11006 34802 11058 34814
rect 7634 34750 7646 34802
rect 7698 34750 7710 34802
rect 5630 34738 5682 34750
rect 11006 34738 11058 34750
rect 11118 34802 11170 34814
rect 18846 34802 18898 34814
rect 33182 34802 33234 34814
rect 39566 34802 39618 34814
rect 11554 34750 11566 34802
rect 11618 34750 11630 34802
rect 14802 34750 14814 34802
rect 14866 34750 14878 34802
rect 15810 34750 15822 34802
rect 15874 34750 15886 34802
rect 16818 34750 16830 34802
rect 16882 34750 16894 34802
rect 21634 34750 21646 34802
rect 21698 34750 21710 34802
rect 24210 34750 24222 34802
rect 24274 34750 24286 34802
rect 25330 34750 25342 34802
rect 25394 34750 25406 34802
rect 26114 34750 26126 34802
rect 26178 34750 26190 34802
rect 34850 34750 34862 34802
rect 34914 34750 34926 34802
rect 36306 34750 36318 34802
rect 36370 34750 36382 34802
rect 37090 34750 37102 34802
rect 37154 34750 37166 34802
rect 11118 34738 11170 34750
rect 18846 34738 18898 34750
rect 33182 34738 33234 34750
rect 39566 34738 39618 34750
rect 1822 34690 1874 34702
rect 1822 34626 1874 34638
rect 2494 34690 2546 34702
rect 2494 34626 2546 34638
rect 6190 34690 6242 34702
rect 6190 34626 6242 34638
rect 12014 34690 12066 34702
rect 12014 34626 12066 34638
rect 12910 34690 12962 34702
rect 19070 34690 19122 34702
rect 13570 34638 13582 34690
rect 13634 34638 13646 34690
rect 13794 34638 13806 34690
rect 13858 34638 13870 34690
rect 12910 34626 12962 34638
rect 19070 34626 19122 34638
rect 19294 34690 19346 34702
rect 19294 34626 19346 34638
rect 20190 34690 20242 34702
rect 20190 34626 20242 34638
rect 20414 34690 20466 34702
rect 28030 34690 28082 34702
rect 22754 34638 22766 34690
rect 22818 34638 22830 34690
rect 20414 34626 20466 34638
rect 28030 34626 28082 34638
rect 28702 34690 28754 34702
rect 28702 34626 28754 34638
rect 32622 34690 32674 34702
rect 35298 34638 35310 34690
rect 35362 34638 35374 34690
rect 37202 34638 37214 34690
rect 37266 34638 37278 34690
rect 32622 34626 32674 34638
rect 1344 34522 58576 34556
rect 1344 34470 19838 34522
rect 19890 34470 19942 34522
rect 19994 34470 20046 34522
rect 20098 34470 50558 34522
rect 50610 34470 50662 34522
rect 50714 34470 50766 34522
rect 50818 34470 58576 34522
rect 1344 34436 58576 34470
rect 1710 34354 1762 34366
rect 1710 34290 1762 34302
rect 3838 34354 3890 34366
rect 3838 34290 3890 34302
rect 5406 34354 5458 34366
rect 5406 34290 5458 34302
rect 6638 34354 6690 34366
rect 6638 34290 6690 34302
rect 7870 34354 7922 34366
rect 7870 34290 7922 34302
rect 11566 34354 11618 34366
rect 18510 34354 18562 34366
rect 23998 34354 24050 34366
rect 13010 34302 13022 34354
rect 13074 34302 13086 34354
rect 13906 34302 13918 34354
rect 13970 34302 13982 34354
rect 15810 34302 15822 34354
rect 15874 34302 15886 34354
rect 21522 34302 21534 34354
rect 21586 34302 21598 34354
rect 11566 34290 11618 34302
rect 18510 34290 18562 34302
rect 23998 34290 24050 34302
rect 24670 34354 24722 34366
rect 24670 34290 24722 34302
rect 29262 34354 29314 34366
rect 29262 34290 29314 34302
rect 29710 34354 29762 34366
rect 29710 34290 29762 34302
rect 30718 34354 30770 34366
rect 30718 34290 30770 34302
rect 10558 34242 10610 34254
rect 15934 34242 15986 34254
rect 2034 34190 2046 34242
rect 2098 34190 2110 34242
rect 14242 34190 14254 34242
rect 14306 34190 14318 34242
rect 14690 34190 14702 34242
rect 14754 34190 14766 34242
rect 10558 34178 10610 34190
rect 15934 34178 15986 34190
rect 17502 34242 17554 34254
rect 17502 34178 17554 34190
rect 18062 34242 18114 34254
rect 28030 34242 28082 34254
rect 19954 34190 19966 34242
rect 20018 34190 20030 34242
rect 21970 34190 21982 34242
rect 22034 34190 22046 34242
rect 23874 34190 23886 34242
rect 23938 34190 23950 34242
rect 18062 34178 18114 34190
rect 28030 34178 28082 34190
rect 28254 34242 28306 34254
rect 28254 34178 28306 34190
rect 35646 34242 35698 34254
rect 35646 34178 35698 34190
rect 8542 34130 8594 34142
rect 10334 34130 10386 34142
rect 9650 34078 9662 34130
rect 9714 34078 9726 34130
rect 8542 34066 8594 34078
rect 10334 34066 10386 34078
rect 10670 34130 10722 34142
rect 10670 34066 10722 34078
rect 12462 34130 12514 34142
rect 16718 34130 16770 34142
rect 12898 34078 12910 34130
rect 12962 34078 12974 34130
rect 14354 34078 14366 34130
rect 14418 34078 14430 34130
rect 15250 34078 15262 34130
rect 15314 34078 15326 34130
rect 16146 34078 16158 34130
rect 16210 34078 16222 34130
rect 12462 34066 12514 34078
rect 16718 34066 16770 34078
rect 17614 34130 17666 34142
rect 17614 34066 17666 34078
rect 18398 34130 18450 34142
rect 18398 34066 18450 34078
rect 18622 34130 18674 34142
rect 18622 34066 18674 34078
rect 19070 34130 19122 34142
rect 19070 34066 19122 34078
rect 19518 34130 19570 34142
rect 22206 34130 22258 34142
rect 28142 34130 28194 34142
rect 36094 34130 36146 34142
rect 20290 34078 20302 34130
rect 20354 34078 20366 34130
rect 20962 34078 20974 34130
rect 21026 34078 21038 34130
rect 21186 34078 21198 34130
rect 21250 34078 21262 34130
rect 22642 34078 22654 34130
rect 22706 34078 22718 34130
rect 23538 34078 23550 34130
rect 23602 34078 23614 34130
rect 23986 34078 23998 34130
rect 24050 34078 24062 34130
rect 25330 34078 25342 34130
rect 25394 34078 25406 34130
rect 25554 34078 25566 34130
rect 25618 34078 25630 34130
rect 26226 34078 26238 34130
rect 26290 34078 26302 34130
rect 33058 34078 33070 34130
rect 33122 34078 33134 34130
rect 19518 34066 19570 34078
rect 22206 34066 22258 34078
rect 28142 34066 28194 34078
rect 36094 34066 36146 34078
rect 36430 34130 36482 34142
rect 39442 34078 39454 34130
rect 39506 34078 39518 34130
rect 36430 34066 36482 34078
rect 2494 34018 2546 34030
rect 7086 34018 7138 34030
rect 3378 33966 3390 34018
rect 3442 33966 3454 34018
rect 5842 33966 5854 34018
rect 5906 33966 5918 34018
rect 2494 33954 2546 33966
rect 7086 33954 7138 33966
rect 7310 34018 7362 34030
rect 7310 33954 7362 33966
rect 8318 34018 8370 34030
rect 8318 33954 8370 33966
rect 10110 34018 10162 34030
rect 10110 33954 10162 33966
rect 11118 34018 11170 34030
rect 27246 34018 27298 34030
rect 12002 33966 12014 34018
rect 12066 33966 12078 34018
rect 11118 33954 11170 33966
rect 27246 33954 27298 33966
rect 28814 34018 28866 34030
rect 36542 34018 36594 34030
rect 30258 33966 30270 34018
rect 30322 33966 30334 34018
rect 34178 33966 34190 34018
rect 34242 33966 34254 34018
rect 38882 33966 38894 34018
rect 38946 33966 38958 34018
rect 28814 33954 28866 33966
rect 36542 33954 36594 33966
rect 8878 33906 8930 33918
rect 8878 33842 8930 33854
rect 17502 33906 17554 33918
rect 17502 33842 17554 33854
rect 26126 33906 26178 33918
rect 27570 33854 27582 33906
rect 27634 33854 27646 33906
rect 26126 33842 26178 33854
rect 1344 33738 58576 33772
rect 1344 33686 4478 33738
rect 4530 33686 4582 33738
rect 4634 33686 4686 33738
rect 4738 33686 35198 33738
rect 35250 33686 35302 33738
rect 35354 33686 35406 33738
rect 35458 33686 58576 33738
rect 1344 33652 58576 33686
rect 18958 33570 19010 33582
rect 14354 33518 14366 33570
rect 14418 33567 14430 33570
rect 14914 33567 14926 33570
rect 14418 33521 14926 33567
rect 14418 33518 14430 33521
rect 14914 33518 14926 33521
rect 14978 33518 14990 33570
rect 16146 33518 16158 33570
rect 16210 33567 16222 33570
rect 16370 33567 16382 33570
rect 16210 33521 16382 33567
rect 16210 33518 16222 33521
rect 16370 33518 16382 33521
rect 16434 33518 16446 33570
rect 18958 33506 19010 33518
rect 32174 33570 32226 33582
rect 32174 33506 32226 33518
rect 9662 33458 9714 33470
rect 7746 33406 7758 33458
rect 7810 33406 7822 33458
rect 9662 33394 9714 33406
rect 14590 33458 14642 33470
rect 14590 33394 14642 33406
rect 15486 33458 15538 33470
rect 20302 33458 20354 33470
rect 17154 33406 17166 33458
rect 17218 33406 17230 33458
rect 15486 33394 15538 33406
rect 20302 33394 20354 33406
rect 23326 33458 23378 33470
rect 27918 33458 27970 33470
rect 26562 33406 26574 33458
rect 26626 33406 26638 33458
rect 23326 33394 23378 33406
rect 27918 33394 27970 33406
rect 2606 33346 2658 33358
rect 2606 33282 2658 33294
rect 3838 33346 3890 33358
rect 3838 33282 3890 33294
rect 4398 33346 4450 33358
rect 4398 33282 4450 33294
rect 4622 33346 4674 33358
rect 19070 33346 19122 33358
rect 27806 33346 27858 33358
rect 5058 33294 5070 33346
rect 5122 33294 5134 33346
rect 5954 33294 5966 33346
rect 6018 33294 6030 33346
rect 9202 33294 9214 33346
rect 9266 33294 9278 33346
rect 17490 33294 17502 33346
rect 17554 33294 17566 33346
rect 18386 33294 18398 33346
rect 18450 33294 18462 33346
rect 23762 33294 23774 33346
rect 23826 33294 23838 33346
rect 25666 33294 25678 33346
rect 25730 33294 25742 33346
rect 4622 33282 4674 33294
rect 19070 33282 19122 33294
rect 27806 33282 27858 33294
rect 28030 33346 28082 33358
rect 28030 33282 28082 33294
rect 30270 33346 30322 33358
rect 35198 33346 35250 33358
rect 37102 33346 37154 33358
rect 41246 33346 41298 33358
rect 30706 33294 30718 33346
rect 30770 33294 30782 33346
rect 33394 33294 33406 33346
rect 33458 33294 33470 33346
rect 36194 33294 36206 33346
rect 36258 33294 36270 33346
rect 39106 33294 39118 33346
rect 39170 33294 39182 33346
rect 30270 33282 30322 33294
rect 35198 33282 35250 33294
rect 37102 33282 37154 33294
rect 41246 33282 41298 33294
rect 1710 33234 1762 33246
rect 1710 33170 1762 33182
rect 3166 33234 3218 33246
rect 3166 33170 3218 33182
rect 3502 33234 3554 33246
rect 3502 33170 3554 33182
rect 4510 33234 4562 33246
rect 18286 33234 18338 33246
rect 28254 33234 28306 33246
rect 7410 33182 7422 33234
rect 7474 33182 7486 33234
rect 8418 33182 8430 33234
rect 8482 33182 8494 33234
rect 17154 33182 17166 33234
rect 17218 33182 17230 33234
rect 25218 33182 25230 33234
rect 25282 33182 25294 33234
rect 26450 33182 26462 33234
rect 26514 33182 26526 33234
rect 4510 33170 4562 33182
rect 18286 33170 18338 33182
rect 28254 33170 28306 33182
rect 29262 33234 29314 33246
rect 38670 33234 38722 33246
rect 32946 33182 32958 33234
rect 33010 33182 33022 33234
rect 33842 33182 33854 33234
rect 33906 33182 33918 33234
rect 29262 33170 29314 33182
rect 38670 33170 38722 33182
rect 40126 33234 40178 33246
rect 40126 33170 40178 33182
rect 2046 33122 2098 33134
rect 2046 33058 2098 33070
rect 3614 33122 3666 33134
rect 3614 33058 3666 33070
rect 10110 33122 10162 33134
rect 10110 33058 10162 33070
rect 12126 33122 12178 33134
rect 12126 33058 12178 33070
rect 12462 33122 12514 33134
rect 12462 33058 12514 33070
rect 13022 33122 13074 33134
rect 13022 33058 13074 33070
rect 13694 33122 13746 33134
rect 13694 33058 13746 33070
rect 14142 33122 14194 33134
rect 14142 33058 14194 33070
rect 15038 33122 15090 33134
rect 15038 33058 15090 33070
rect 16382 33122 16434 33134
rect 16382 33058 16434 33070
rect 18958 33122 19010 33134
rect 18958 33058 19010 33070
rect 19518 33122 19570 33134
rect 19518 33058 19570 33070
rect 20750 33122 20802 33134
rect 20750 33058 20802 33070
rect 21646 33122 21698 33134
rect 21646 33058 21698 33070
rect 22094 33122 22146 33134
rect 22094 33058 22146 33070
rect 22542 33122 22594 33134
rect 22542 33058 22594 33070
rect 22990 33122 23042 33134
rect 22990 33058 23042 33070
rect 23214 33122 23266 33134
rect 23214 33058 23266 33070
rect 23438 33122 23490 33134
rect 23438 33058 23490 33070
rect 27694 33122 27746 33134
rect 37214 33122 37266 33134
rect 36418 33070 36430 33122
rect 36482 33070 36494 33122
rect 37650 33070 37662 33122
rect 37714 33070 37726 33122
rect 27694 33058 27746 33070
rect 37214 33058 37266 33070
rect 1344 32954 58576 32988
rect 1344 32902 19838 32954
rect 19890 32902 19942 32954
rect 19994 32902 20046 32954
rect 20098 32902 50558 32954
rect 50610 32902 50662 32954
rect 50714 32902 50766 32954
rect 50818 32902 58576 32954
rect 1344 32868 58576 32902
rect 19182 32786 19234 32798
rect 6738 32734 6750 32786
rect 6802 32734 6814 32786
rect 13458 32734 13470 32786
rect 13522 32734 13534 32786
rect 19182 32722 19234 32734
rect 28926 32786 28978 32798
rect 40910 32786 40962 32798
rect 34066 32734 34078 32786
rect 34130 32734 34142 32786
rect 28926 32722 28978 32734
rect 40910 32722 40962 32734
rect 13918 32674 13970 32686
rect 5394 32622 5406 32674
rect 5458 32622 5470 32674
rect 13918 32610 13970 32622
rect 14254 32674 14306 32686
rect 28366 32674 28418 32686
rect 18050 32622 18062 32674
rect 18114 32622 18126 32674
rect 21858 32622 21870 32674
rect 21922 32622 21934 32674
rect 22306 32622 22318 32674
rect 22370 32622 22382 32674
rect 22754 32622 22766 32674
rect 22818 32622 22830 32674
rect 14254 32610 14306 32622
rect 28366 32610 28418 32622
rect 28478 32674 28530 32686
rect 35646 32674 35698 32686
rect 41470 32674 41522 32686
rect 33170 32622 33182 32674
rect 33234 32622 33246 32674
rect 37314 32622 37326 32674
rect 37378 32622 37390 32674
rect 28478 32610 28530 32622
rect 35646 32610 35698 32622
rect 41470 32610 41522 32622
rect 7310 32562 7362 32574
rect 2930 32510 2942 32562
rect 2994 32510 3006 32562
rect 3266 32510 3278 32562
rect 3330 32510 3342 32562
rect 3602 32510 3614 32562
rect 3666 32510 3678 32562
rect 4946 32510 4958 32562
rect 5010 32510 5022 32562
rect 6514 32510 6526 32562
rect 6578 32510 6590 32562
rect 7310 32498 7362 32510
rect 8990 32562 9042 32574
rect 13134 32562 13186 32574
rect 10434 32510 10446 32562
rect 10498 32510 10510 32562
rect 12786 32510 12798 32562
rect 12850 32510 12862 32562
rect 8990 32498 9042 32510
rect 13134 32498 13186 32510
rect 16830 32562 16882 32574
rect 28142 32562 28194 32574
rect 35198 32562 35250 32574
rect 17714 32510 17726 32562
rect 17778 32510 17790 32562
rect 18834 32510 18846 32562
rect 18898 32510 18910 32562
rect 21634 32510 21646 32562
rect 21698 32510 21710 32562
rect 23650 32510 23662 32562
rect 23714 32510 23726 32562
rect 25330 32510 25342 32562
rect 25394 32510 25406 32562
rect 27682 32510 27694 32562
rect 27746 32510 27758 32562
rect 34626 32510 34638 32562
rect 34690 32510 34702 32562
rect 38434 32510 38446 32562
rect 38498 32510 38510 32562
rect 38770 32510 38782 32562
rect 38834 32510 38846 32562
rect 16830 32498 16882 32510
rect 28142 32498 28194 32510
rect 35198 32498 35250 32510
rect 15262 32450 15314 32462
rect 8530 32398 8542 32450
rect 8594 32398 8606 32450
rect 10658 32398 10670 32450
rect 10722 32398 10734 32450
rect 14690 32398 14702 32450
rect 14754 32398 14766 32450
rect 15262 32386 15314 32398
rect 16494 32450 16546 32462
rect 19854 32450 19906 32462
rect 18050 32398 18062 32450
rect 18114 32398 18126 32450
rect 16494 32386 16546 32398
rect 19854 32386 19906 32398
rect 21422 32450 21474 32462
rect 21422 32386 21474 32398
rect 24670 32450 24722 32462
rect 27794 32398 27806 32450
rect 27858 32398 27870 32450
rect 39442 32398 39454 32450
rect 39506 32398 39518 32450
rect 24670 32386 24722 32398
rect 10770 32286 10782 32338
rect 10834 32286 10846 32338
rect 26786 32286 26798 32338
rect 26850 32286 26862 32338
rect 1344 32170 58576 32204
rect 1344 32118 4478 32170
rect 4530 32118 4582 32170
rect 4634 32118 4686 32170
rect 4738 32118 35198 32170
rect 35250 32118 35302 32170
rect 35354 32118 35406 32170
rect 35458 32118 58576 32170
rect 1344 32084 58576 32118
rect 17054 32002 17106 32014
rect 17054 31938 17106 31950
rect 25006 32002 25058 32014
rect 25006 31938 25058 31950
rect 3726 31890 3778 31902
rect 20862 31890 20914 31902
rect 2930 31838 2942 31890
rect 2994 31838 3006 31890
rect 15138 31838 15150 31890
rect 15202 31838 15214 31890
rect 3726 31826 3778 31838
rect 20862 31826 20914 31838
rect 23438 31890 23490 31902
rect 23438 31826 23490 31838
rect 27134 31890 27186 31902
rect 27134 31826 27186 31838
rect 29150 31890 29202 31902
rect 29150 31826 29202 31838
rect 30382 31890 30434 31902
rect 30382 31826 30434 31838
rect 33854 31890 33906 31902
rect 33854 31826 33906 31838
rect 4286 31778 4338 31790
rect 13470 31778 13522 31790
rect 3266 31726 3278 31778
rect 3330 31726 3342 31778
rect 8978 31726 8990 31778
rect 9042 31726 9054 31778
rect 9314 31726 9326 31778
rect 9378 31726 9390 31778
rect 9650 31726 9662 31778
rect 9714 31726 9726 31778
rect 10994 31726 11006 31778
rect 11058 31726 11070 31778
rect 12786 31726 12798 31778
rect 12850 31726 12862 31778
rect 4286 31714 4338 31726
rect 13470 31714 13522 31726
rect 14030 31778 14082 31790
rect 14030 31714 14082 31726
rect 14814 31778 14866 31790
rect 14814 31714 14866 31726
rect 15038 31778 15090 31790
rect 20078 31778 20130 31790
rect 15810 31726 15822 31778
rect 15874 31726 15886 31778
rect 16594 31726 16606 31778
rect 16658 31726 16670 31778
rect 17042 31726 17054 31778
rect 17106 31726 17118 31778
rect 17602 31726 17614 31778
rect 17666 31726 17678 31778
rect 18498 31726 18510 31778
rect 18562 31726 18574 31778
rect 19506 31726 19518 31778
rect 19570 31726 19582 31778
rect 15038 31714 15090 31726
rect 20078 31714 20130 31726
rect 20190 31778 20242 31790
rect 20190 31714 20242 31726
rect 20526 31778 20578 31790
rect 20526 31714 20578 31726
rect 22318 31778 22370 31790
rect 26798 31778 26850 31790
rect 33742 31778 33794 31790
rect 22754 31726 22766 31778
rect 22818 31726 22830 31778
rect 24994 31726 25006 31778
rect 25058 31726 25070 31778
rect 28242 31726 28254 31778
rect 28306 31726 28318 31778
rect 22318 31714 22370 31726
rect 26798 31714 26850 31726
rect 33742 31714 33794 31726
rect 34190 31778 34242 31790
rect 34190 31714 34242 31726
rect 38670 31778 38722 31790
rect 38670 31714 38722 31726
rect 39118 31778 39170 31790
rect 39118 31714 39170 31726
rect 11902 31666 11954 31678
rect 11902 31602 11954 31614
rect 14590 31666 14642 31678
rect 14590 31602 14642 31614
rect 16046 31666 16098 31678
rect 21422 31666 21474 31678
rect 33182 31666 33234 31678
rect 17714 31614 17726 31666
rect 17778 31614 17790 31666
rect 24210 31614 24222 31666
rect 24274 31614 24286 31666
rect 25218 31614 25230 31666
rect 25282 31614 25294 31666
rect 27794 31614 27806 31666
rect 27858 31614 27870 31666
rect 28018 31614 28030 31666
rect 28082 31614 28094 31666
rect 16046 31602 16098 31614
rect 21422 31602 21474 31614
rect 33182 31602 33234 31614
rect 35198 31666 35250 31678
rect 39678 31666 39730 31678
rect 36978 31614 36990 31666
rect 37042 31614 37054 31666
rect 35198 31602 35250 31614
rect 39678 31602 39730 31614
rect 15150 31554 15202 31566
rect 19742 31554 19794 31566
rect 12898 31502 12910 31554
rect 12962 31502 12974 31554
rect 18050 31502 18062 31554
rect 18114 31502 18126 31554
rect 18946 31502 18958 31554
rect 19010 31502 19022 31554
rect 15150 31490 15202 31502
rect 19742 31490 19794 31502
rect 20302 31554 20354 31566
rect 20302 31490 20354 31502
rect 29710 31554 29762 31566
rect 29710 31490 29762 31502
rect 30942 31554 30994 31566
rect 37202 31502 37214 31554
rect 37266 31502 37278 31554
rect 30942 31490 30994 31502
rect 1344 31386 58576 31420
rect 1344 31334 19838 31386
rect 19890 31334 19942 31386
rect 19994 31334 20046 31386
rect 20098 31334 50558 31386
rect 50610 31334 50662 31386
rect 50714 31334 50766 31386
rect 50818 31334 58576 31386
rect 1344 31300 58576 31334
rect 2270 31218 2322 31230
rect 2270 31154 2322 31166
rect 7534 31218 7586 31230
rect 7534 31154 7586 31166
rect 9102 31218 9154 31230
rect 14142 31218 14194 31230
rect 10882 31166 10894 31218
rect 10946 31166 10958 31218
rect 13122 31166 13134 31218
rect 13186 31166 13198 31218
rect 9102 31154 9154 31166
rect 14142 31154 14194 31166
rect 15150 31218 15202 31230
rect 15150 31154 15202 31166
rect 16270 31218 16322 31230
rect 16270 31154 16322 31166
rect 17838 31218 17890 31230
rect 18734 31218 18786 31230
rect 18050 31166 18062 31218
rect 18114 31166 18126 31218
rect 17838 31154 17890 31166
rect 18734 31154 18786 31166
rect 19070 31218 19122 31230
rect 19070 31154 19122 31166
rect 20974 31218 21026 31230
rect 20974 31154 21026 31166
rect 23886 31218 23938 31230
rect 23886 31154 23938 31166
rect 25790 31218 25842 31230
rect 25790 31154 25842 31166
rect 26126 31218 26178 31230
rect 26126 31154 26178 31166
rect 26350 31218 26402 31230
rect 26350 31154 26402 31166
rect 26574 31218 26626 31230
rect 26574 31154 26626 31166
rect 27582 31218 27634 31230
rect 27582 31154 27634 31166
rect 27806 31218 27858 31230
rect 27806 31154 27858 31166
rect 27918 31218 27970 31230
rect 27918 31154 27970 31166
rect 28926 31218 28978 31230
rect 33170 31166 33182 31218
rect 33234 31166 33246 31218
rect 28926 31154 28978 31166
rect 13918 31106 13970 31118
rect 3042 31054 3054 31106
rect 3106 31054 3118 31106
rect 4386 31054 4398 31106
rect 4450 31054 4462 31106
rect 5618 31054 5630 31106
rect 5682 31054 5694 31106
rect 12562 31054 12574 31106
rect 12626 31054 12638 31106
rect 13918 31042 13970 31054
rect 15486 31106 15538 31118
rect 15486 31042 15538 31054
rect 17390 31106 17442 31118
rect 17390 31042 17442 31054
rect 17614 31106 17666 31118
rect 17614 31042 17666 31054
rect 18510 31106 18562 31118
rect 18510 31042 18562 31054
rect 18846 31106 18898 31118
rect 18846 31042 18898 31054
rect 20078 31106 20130 31118
rect 20078 31042 20130 31054
rect 20302 31106 20354 31118
rect 24446 31106 24498 31118
rect 21074 31054 21086 31106
rect 21138 31103 21150 31106
rect 21298 31103 21310 31106
rect 21138 31057 21310 31103
rect 21138 31054 21150 31057
rect 21298 31054 21310 31057
rect 21362 31054 21374 31106
rect 20302 31042 20354 31054
rect 24446 31042 24498 31054
rect 24670 31106 24722 31118
rect 24670 31042 24722 31054
rect 34302 31106 34354 31118
rect 34302 31042 34354 31054
rect 35758 31106 35810 31118
rect 35758 31042 35810 31054
rect 14366 30994 14418 31006
rect 16158 30994 16210 31006
rect 2034 30942 2046 30994
rect 2098 30942 2110 30994
rect 3490 30942 3502 30994
rect 3554 30942 3566 30994
rect 4834 30942 4846 30994
rect 4898 30942 4910 30994
rect 5506 30942 5518 30994
rect 5570 30942 5582 30994
rect 10098 30942 10110 30994
rect 10162 30942 10174 30994
rect 10994 30942 11006 30994
rect 11058 30942 11070 30994
rect 11778 30942 11790 30994
rect 11842 30942 11854 30994
rect 13346 30942 13358 30994
rect 13410 30942 13422 30994
rect 14578 30942 14590 30994
rect 14642 30942 14654 30994
rect 14366 30930 14418 30942
rect 16158 30930 16210 30942
rect 16830 30994 16882 31006
rect 16830 30930 16882 30942
rect 18062 30994 18114 31006
rect 18062 30930 18114 30942
rect 18958 30994 19010 31006
rect 18958 30930 19010 30942
rect 20638 30994 20690 31006
rect 26238 30994 26290 31006
rect 24210 30942 24222 30994
rect 24274 30942 24286 30994
rect 20638 30930 20690 30942
rect 26238 30930 26290 30942
rect 28030 30994 28082 31006
rect 28030 30930 28082 30942
rect 28702 30994 28754 31006
rect 28702 30930 28754 30942
rect 29374 30994 29426 31006
rect 29374 30930 29426 30942
rect 34750 30994 34802 31006
rect 36866 30942 36878 30994
rect 36930 30942 36942 30994
rect 38210 30942 38222 30994
rect 38274 30942 38286 30994
rect 34750 30930 34802 30942
rect 8654 30882 8706 30894
rect 3378 30830 3390 30882
rect 3442 30830 3454 30882
rect 6290 30830 6302 30882
rect 6354 30830 6366 30882
rect 8654 30818 8706 30830
rect 14254 30882 14306 30894
rect 14254 30818 14306 30830
rect 19630 30882 19682 30894
rect 19630 30818 19682 30830
rect 21422 30882 21474 30894
rect 21422 30818 21474 30830
rect 21870 30882 21922 30894
rect 27134 30882 27186 30894
rect 28814 30882 28866 30894
rect 24546 30830 24558 30882
rect 24610 30830 24622 30882
rect 25330 30830 25342 30882
rect 25394 30830 25406 30882
rect 27458 30879 27470 30882
rect 21870 30818 21922 30830
rect 27134 30818 27186 30830
rect 27249 30833 27470 30879
rect 16270 30770 16322 30782
rect 8642 30718 8654 30770
rect 8706 30767 8718 30770
rect 9090 30767 9102 30770
rect 8706 30721 9102 30767
rect 8706 30718 8718 30721
rect 9090 30718 9102 30721
rect 9154 30718 9166 30770
rect 16270 30706 16322 30718
rect 20862 30770 20914 30782
rect 27249 30770 27295 30833
rect 27458 30830 27470 30833
rect 27522 30830 27534 30882
rect 37426 30830 37438 30882
rect 37490 30830 37502 30882
rect 28814 30818 28866 30830
rect 21074 30718 21086 30770
rect 21138 30767 21150 30770
rect 21858 30767 21870 30770
rect 21138 30721 21870 30767
rect 21138 30718 21150 30721
rect 21858 30718 21870 30721
rect 21922 30718 21934 30770
rect 27234 30718 27246 30770
rect 27298 30718 27310 30770
rect 20862 30706 20914 30718
rect 1344 30602 58576 30636
rect 1344 30550 4478 30602
rect 4530 30550 4582 30602
rect 4634 30550 4686 30602
rect 4738 30550 35198 30602
rect 35250 30550 35302 30602
rect 35354 30550 35406 30602
rect 35458 30550 58576 30602
rect 1344 30516 58576 30550
rect 4958 30434 5010 30446
rect 21422 30434 21474 30446
rect 14354 30382 14366 30434
rect 14418 30431 14430 30434
rect 14690 30431 14702 30434
rect 14418 30385 14702 30431
rect 14418 30382 14430 30385
rect 14690 30382 14702 30385
rect 14754 30382 14766 30434
rect 4958 30370 5010 30382
rect 21422 30370 21474 30382
rect 14702 30322 14754 30334
rect 6626 30270 6638 30322
rect 6690 30270 6702 30322
rect 11554 30270 11566 30322
rect 11618 30270 11630 30322
rect 14702 30258 14754 30270
rect 15262 30322 15314 30334
rect 15262 30258 15314 30270
rect 17166 30322 17218 30334
rect 17166 30258 17218 30270
rect 26350 30322 26402 30334
rect 26350 30258 26402 30270
rect 27134 30322 27186 30334
rect 27134 30258 27186 30270
rect 28366 30322 28418 30334
rect 31502 30322 31554 30334
rect 30482 30270 30494 30322
rect 30546 30270 30558 30322
rect 28366 30258 28418 30270
rect 31502 30258 31554 30270
rect 34526 30322 34578 30334
rect 34526 30258 34578 30270
rect 1710 30210 1762 30222
rect 9102 30210 9154 30222
rect 6850 30158 6862 30210
rect 6914 30158 6926 30210
rect 7858 30158 7870 30210
rect 7922 30158 7934 30210
rect 8642 30158 8654 30210
rect 8706 30158 8718 30210
rect 1710 30146 1762 30158
rect 9102 30146 9154 30158
rect 9886 30210 9938 30222
rect 12910 30210 12962 30222
rect 11442 30158 11454 30210
rect 11506 30158 11518 30210
rect 9886 30146 9938 30158
rect 12910 30146 12962 30158
rect 17502 30210 17554 30222
rect 21534 30210 21586 30222
rect 17714 30158 17726 30210
rect 17778 30158 17790 30210
rect 20066 30158 20078 30210
rect 20130 30158 20142 30210
rect 17502 30146 17554 30158
rect 21534 30146 21586 30158
rect 21758 30210 21810 30222
rect 23550 30210 23602 30222
rect 22530 30158 22542 30210
rect 22594 30158 22606 30210
rect 21758 30146 21810 30158
rect 23550 30146 23602 30158
rect 25118 30210 25170 30222
rect 25118 30146 25170 30158
rect 25230 30210 25282 30222
rect 37214 30210 37266 30222
rect 25554 30158 25566 30210
rect 25618 30158 25630 30210
rect 30930 30158 30942 30210
rect 30994 30158 31006 30210
rect 31938 30158 31950 30210
rect 32002 30158 32014 30210
rect 34962 30158 34974 30210
rect 35026 30158 35038 30210
rect 35634 30158 35646 30210
rect 35698 30158 35710 30210
rect 25230 30146 25282 30158
rect 37214 30146 37266 30158
rect 2046 30098 2098 30110
rect 2046 30034 2098 30046
rect 2382 30098 2434 30110
rect 2382 30034 2434 30046
rect 5070 30098 5122 30110
rect 5070 30034 5122 30046
rect 6190 30098 6242 30110
rect 6190 30034 6242 30046
rect 6638 30098 6690 30110
rect 11678 30098 11730 30110
rect 7522 30046 7534 30098
rect 7586 30046 7598 30098
rect 9650 30046 9662 30098
rect 9714 30046 9726 30098
rect 6638 30034 6690 30046
rect 11678 30034 11730 30046
rect 12126 30098 12178 30110
rect 12126 30034 12178 30046
rect 12574 30098 12626 30110
rect 21310 30098 21362 30110
rect 19954 30046 19966 30098
rect 20018 30046 20030 30098
rect 12574 30034 12626 30046
rect 21310 30034 21362 30046
rect 21982 30098 22034 30110
rect 25342 30098 25394 30110
rect 22642 30046 22654 30098
rect 22706 30046 22718 30098
rect 23202 30046 23214 30098
rect 23266 30046 23278 30098
rect 24098 30046 24110 30098
rect 24162 30046 24174 30098
rect 24546 30046 24558 30098
rect 24610 30046 24622 30098
rect 21982 30034 22034 30046
rect 25342 30034 25394 30046
rect 35982 30098 36034 30110
rect 35982 30034 36034 30046
rect 36542 30098 36594 30110
rect 36542 30034 36594 30046
rect 2718 29986 2770 29998
rect 2718 29922 2770 29934
rect 3166 29986 3218 29998
rect 3166 29922 3218 29934
rect 4174 29986 4226 29998
rect 4174 29922 4226 29934
rect 4622 29986 4674 29998
rect 4622 29922 4674 29934
rect 4958 29986 5010 29998
rect 4958 29922 5010 29934
rect 5854 29986 5906 29998
rect 5854 29922 5906 29934
rect 6414 29986 6466 29998
rect 10670 29986 10722 29998
rect 7746 29934 7758 29986
rect 7810 29934 7822 29986
rect 6414 29922 6466 29934
rect 10670 29922 10722 29934
rect 11230 29986 11282 29998
rect 11230 29922 11282 29934
rect 11902 29986 11954 29998
rect 11902 29922 11954 29934
rect 12686 29986 12738 29998
rect 12686 29922 12738 29934
rect 13582 29986 13634 29998
rect 13582 29922 13634 29934
rect 14254 29986 14306 29998
rect 26014 29986 26066 29998
rect 19170 29934 19182 29986
rect 19234 29934 19246 29986
rect 23986 29934 23998 29986
rect 24050 29934 24062 29986
rect 14254 29922 14306 29934
rect 26014 29922 26066 29934
rect 29262 29986 29314 29998
rect 29262 29922 29314 29934
rect 1344 29818 58576 29852
rect 1344 29766 19838 29818
rect 19890 29766 19942 29818
rect 19994 29766 20046 29818
rect 20098 29766 50558 29818
rect 50610 29766 50662 29818
rect 50714 29766 50766 29818
rect 50818 29766 58576 29818
rect 1344 29732 58576 29766
rect 1822 29650 1874 29662
rect 7086 29650 7138 29662
rect 18958 29650 19010 29662
rect 6178 29598 6190 29650
rect 6242 29598 6254 29650
rect 15138 29598 15150 29650
rect 15202 29598 15214 29650
rect 1822 29586 1874 29598
rect 7086 29586 7138 29598
rect 18958 29586 19010 29598
rect 19518 29650 19570 29662
rect 19518 29586 19570 29598
rect 20078 29650 20130 29662
rect 20078 29586 20130 29598
rect 23550 29650 23602 29662
rect 23550 29586 23602 29598
rect 23886 29650 23938 29662
rect 23886 29586 23938 29598
rect 24110 29650 24162 29662
rect 24110 29586 24162 29598
rect 24334 29650 24386 29662
rect 24334 29586 24386 29598
rect 25902 29650 25954 29662
rect 25902 29586 25954 29598
rect 27134 29650 27186 29662
rect 27134 29586 27186 29598
rect 27694 29650 27746 29662
rect 35746 29598 35758 29650
rect 35810 29598 35822 29650
rect 27694 29586 27746 29598
rect 11790 29538 11842 29550
rect 3154 29486 3166 29538
rect 3218 29486 3230 29538
rect 6402 29486 6414 29538
rect 6466 29486 6478 29538
rect 7410 29486 7422 29538
rect 7474 29486 7486 29538
rect 9762 29486 9774 29538
rect 9826 29486 9838 29538
rect 11790 29474 11842 29486
rect 13694 29538 13746 29550
rect 13694 29474 13746 29486
rect 13918 29538 13970 29550
rect 13918 29474 13970 29486
rect 14702 29538 14754 29550
rect 14702 29474 14754 29486
rect 20414 29538 20466 29550
rect 20414 29474 20466 29486
rect 22430 29538 22482 29550
rect 37438 29538 37490 29550
rect 29586 29486 29598 29538
rect 29650 29486 29662 29538
rect 34290 29486 34302 29538
rect 34354 29486 34366 29538
rect 22430 29474 22482 29486
rect 37438 29474 37490 29486
rect 13358 29426 13410 29438
rect 14590 29426 14642 29438
rect 19966 29426 20018 29438
rect 2258 29374 2270 29426
rect 2322 29374 2334 29426
rect 4610 29374 4622 29426
rect 4674 29374 4686 29426
rect 5730 29374 5742 29426
rect 5794 29374 5806 29426
rect 7522 29374 7534 29426
rect 7586 29374 7598 29426
rect 7970 29374 7982 29426
rect 8034 29374 8046 29426
rect 8866 29374 8878 29426
rect 8930 29374 8942 29426
rect 9650 29374 9662 29426
rect 9714 29374 9726 29426
rect 10210 29374 10222 29426
rect 10274 29374 10286 29426
rect 10994 29374 11006 29426
rect 11058 29374 11070 29426
rect 12450 29374 12462 29426
rect 12514 29374 12526 29426
rect 14354 29374 14366 29426
rect 14418 29374 14430 29426
rect 19730 29374 19742 29426
rect 19794 29374 19806 29426
rect 13358 29362 13410 29374
rect 14590 29362 14642 29374
rect 19966 29362 20018 29374
rect 20190 29426 20242 29438
rect 20190 29362 20242 29374
rect 20974 29426 21026 29438
rect 20974 29362 21026 29374
rect 21534 29426 21586 29438
rect 21534 29362 21586 29374
rect 21982 29426 22034 29438
rect 21982 29362 22034 29374
rect 24446 29426 24498 29438
rect 24446 29362 24498 29374
rect 27246 29426 27298 29438
rect 27246 29362 27298 29374
rect 27918 29426 27970 29438
rect 28354 29374 28366 29426
rect 28418 29374 28430 29426
rect 28802 29374 28814 29426
rect 28866 29374 28878 29426
rect 29474 29374 29486 29426
rect 29538 29374 29550 29426
rect 35858 29374 35870 29426
rect 35922 29374 35934 29426
rect 38098 29374 38110 29426
rect 38162 29374 38174 29426
rect 27918 29362 27970 29374
rect 15598 29314 15650 29326
rect 12114 29262 12126 29314
rect 12178 29262 12190 29314
rect 15598 29250 15650 29262
rect 26574 29314 26626 29326
rect 26574 29250 26626 29262
rect 27806 29314 27858 29326
rect 27806 29250 27858 29262
rect 10222 29202 10274 29214
rect 10222 29138 10274 29150
rect 13134 29202 13186 29214
rect 13134 29138 13186 29150
rect 13806 29202 13858 29214
rect 29026 29150 29038 29202
rect 29090 29150 29102 29202
rect 13806 29138 13858 29150
rect 1344 29034 58576 29068
rect 1344 28982 4478 29034
rect 4530 28982 4582 29034
rect 4634 28982 4686 29034
rect 4738 28982 35198 29034
rect 35250 28982 35302 29034
rect 35354 28982 35406 29034
rect 35458 28982 58576 29034
rect 1344 28948 58576 28982
rect 21422 28866 21474 28878
rect 30146 28814 30158 28866
rect 30210 28814 30222 28866
rect 21422 28802 21474 28814
rect 2606 28754 2658 28766
rect 11902 28754 11954 28766
rect 3826 28702 3838 28754
rect 3890 28702 3902 28754
rect 10770 28702 10782 28754
rect 10834 28702 10846 28754
rect 2606 28690 2658 28702
rect 11902 28690 11954 28702
rect 12238 28754 12290 28766
rect 12238 28690 12290 28702
rect 12686 28754 12738 28766
rect 12686 28690 12738 28702
rect 15038 28754 15090 28766
rect 15038 28690 15090 28702
rect 16718 28754 16770 28766
rect 16718 28690 16770 28702
rect 18174 28754 18226 28766
rect 18174 28690 18226 28702
rect 19182 28754 19234 28766
rect 19182 28690 19234 28702
rect 20078 28754 20130 28766
rect 26910 28754 26962 28766
rect 26338 28702 26350 28754
rect 26402 28702 26414 28754
rect 20078 28690 20130 28702
rect 26910 28690 26962 28702
rect 27358 28754 27410 28766
rect 27358 28690 27410 28702
rect 2382 28642 2434 28654
rect 2382 28578 2434 28590
rect 2830 28642 2882 28654
rect 6190 28642 6242 28654
rect 10222 28642 10274 28654
rect 14478 28642 14530 28654
rect 3938 28590 3950 28642
rect 4002 28590 4014 28642
rect 6514 28590 6526 28642
rect 6578 28590 6590 28642
rect 11330 28590 11342 28642
rect 11394 28590 11406 28642
rect 2830 28578 2882 28590
rect 6190 28578 6242 28590
rect 10222 28578 10274 28590
rect 14478 28578 14530 28590
rect 15262 28642 15314 28654
rect 15262 28578 15314 28590
rect 15822 28642 15874 28654
rect 15822 28578 15874 28590
rect 16158 28642 16210 28654
rect 16158 28578 16210 28590
rect 18734 28642 18786 28654
rect 18734 28578 18786 28590
rect 20414 28642 20466 28654
rect 20414 28578 20466 28590
rect 20750 28642 20802 28654
rect 20750 28578 20802 28590
rect 21870 28642 21922 28654
rect 22878 28642 22930 28654
rect 25118 28642 25170 28654
rect 28478 28642 28530 28654
rect 22306 28590 22318 28642
rect 22370 28590 22382 28642
rect 23538 28590 23550 28642
rect 23602 28590 23614 28642
rect 24098 28590 24110 28642
rect 24162 28590 24174 28642
rect 26002 28590 26014 28642
rect 26066 28590 26078 28642
rect 21870 28578 21922 28590
rect 22878 28578 22930 28590
rect 25118 28578 25170 28590
rect 28478 28578 28530 28590
rect 29150 28642 29202 28654
rect 29150 28578 29202 28590
rect 29262 28642 29314 28654
rect 29262 28578 29314 28590
rect 29598 28642 29650 28654
rect 29598 28578 29650 28590
rect 29710 28642 29762 28654
rect 29710 28578 29762 28590
rect 3278 28530 3330 28542
rect 3278 28466 3330 28478
rect 7086 28530 7138 28542
rect 11118 28530 11170 28542
rect 10322 28478 10334 28530
rect 10386 28478 10398 28530
rect 7086 28466 7138 28478
rect 11118 28466 11170 28478
rect 14702 28530 14754 28542
rect 14702 28466 14754 28478
rect 14926 28530 14978 28542
rect 14926 28466 14978 28478
rect 18622 28530 18674 28542
rect 18622 28466 18674 28478
rect 21534 28530 21586 28542
rect 21534 28466 21586 28478
rect 23438 28530 23490 28542
rect 28142 28530 28194 28542
rect 24210 28478 24222 28530
rect 24274 28478 24286 28530
rect 23438 28466 23490 28478
rect 28142 28466 28194 28478
rect 28254 28530 28306 28542
rect 28254 28466 28306 28478
rect 2494 28418 2546 28430
rect 2494 28354 2546 28366
rect 2718 28418 2770 28430
rect 2718 28354 2770 28366
rect 3502 28418 3554 28430
rect 3502 28354 3554 28366
rect 3726 28418 3778 28430
rect 3726 28354 3778 28366
rect 4398 28418 4450 28430
rect 10782 28418 10834 28430
rect 7970 28366 7982 28418
rect 8034 28366 8046 28418
rect 4398 28354 4450 28366
rect 10782 28354 10834 28366
rect 10894 28418 10946 28430
rect 10894 28354 10946 28366
rect 15150 28418 15202 28430
rect 15150 28354 15202 28366
rect 18398 28418 18450 28430
rect 18398 28354 18450 28366
rect 20526 28418 20578 28430
rect 20526 28354 20578 28366
rect 21422 28418 21474 28430
rect 27918 28418 27970 28430
rect 24322 28366 24334 28418
rect 24386 28366 24398 28418
rect 21422 28354 21474 28366
rect 27918 28354 27970 28366
rect 1344 28250 58576 28284
rect 1344 28198 19838 28250
rect 19890 28198 19942 28250
rect 19994 28198 20046 28250
rect 20098 28198 50558 28250
rect 50610 28198 50662 28250
rect 50714 28198 50766 28250
rect 50818 28198 58576 28250
rect 1344 28164 58576 28198
rect 2046 28082 2098 28094
rect 2046 28018 2098 28030
rect 3950 28082 4002 28094
rect 3950 28018 4002 28030
rect 4846 28082 4898 28094
rect 4846 28018 4898 28030
rect 5294 28082 5346 28094
rect 5294 28018 5346 28030
rect 7198 28082 7250 28094
rect 7198 28018 7250 28030
rect 8542 28082 8594 28094
rect 8542 28018 8594 28030
rect 8654 28082 8706 28094
rect 8654 28018 8706 28030
rect 8766 28082 8818 28094
rect 8766 28018 8818 28030
rect 11566 28082 11618 28094
rect 18174 28082 18226 28094
rect 25342 28082 25394 28094
rect 13010 28030 13022 28082
rect 13074 28030 13086 28082
rect 18386 28030 18398 28082
rect 18450 28030 18462 28082
rect 11566 28018 11618 28030
rect 18174 28018 18226 28030
rect 25342 28018 25394 28030
rect 25678 28082 25730 28094
rect 29710 28082 29762 28094
rect 27010 28030 27022 28082
rect 27074 28030 27086 28082
rect 25678 28018 25730 28030
rect 29710 28018 29762 28030
rect 30606 28082 30658 28094
rect 30606 28018 30658 28030
rect 3726 27970 3778 27982
rect 3726 27906 3778 27918
rect 5070 27970 5122 27982
rect 5070 27906 5122 27918
rect 6078 27970 6130 27982
rect 8990 27970 9042 27982
rect 16718 27970 16770 27982
rect 21646 27970 21698 27982
rect 7970 27918 7982 27970
rect 8034 27918 8046 27970
rect 12338 27918 12350 27970
rect 12402 27918 12414 27970
rect 20514 27918 20526 27970
rect 20578 27918 20590 27970
rect 20962 27918 20974 27970
rect 21026 27918 21038 27970
rect 27346 27918 27358 27970
rect 27410 27918 27422 27970
rect 6078 27906 6130 27918
rect 8990 27906 9042 27918
rect 16718 27906 16770 27918
rect 21646 27906 21698 27918
rect 1710 27858 1762 27870
rect 1710 27794 1762 27806
rect 4286 27858 4338 27870
rect 8430 27858 8482 27870
rect 15710 27858 15762 27870
rect 5506 27806 5518 27858
rect 5570 27806 5582 27858
rect 5842 27806 5854 27858
rect 5906 27806 5918 27858
rect 6738 27806 6750 27858
rect 6802 27806 6814 27858
rect 7074 27806 7086 27858
rect 7138 27806 7150 27858
rect 7746 27806 7758 27858
rect 7810 27806 7822 27858
rect 10770 27806 10782 27858
rect 10834 27806 10846 27858
rect 12114 27806 12126 27858
rect 12178 27806 12190 27858
rect 13682 27806 13694 27858
rect 13746 27806 13758 27858
rect 14242 27806 14254 27858
rect 14306 27806 14318 27858
rect 15474 27806 15486 27858
rect 15538 27806 15550 27858
rect 4286 27794 4338 27806
rect 8430 27794 8482 27806
rect 15710 27794 15762 27806
rect 15822 27858 15874 27870
rect 15822 27794 15874 27806
rect 16606 27858 16658 27870
rect 16606 27794 16658 27806
rect 17726 27858 17778 27870
rect 17726 27794 17778 27806
rect 17950 27858 18002 27870
rect 17950 27794 18002 27806
rect 18398 27858 18450 27870
rect 25230 27858 25282 27870
rect 18722 27806 18734 27858
rect 18786 27806 18798 27858
rect 19394 27806 19406 27858
rect 19458 27806 19470 27858
rect 19954 27806 19966 27858
rect 20018 27806 20030 27858
rect 20402 27806 20414 27858
rect 20466 27806 20478 27858
rect 18398 27794 18450 27806
rect 25230 27794 25282 27806
rect 25454 27858 25506 27870
rect 25454 27794 25506 27806
rect 26462 27858 26514 27870
rect 26462 27794 26514 27806
rect 26686 27858 26738 27870
rect 30046 27858 30098 27870
rect 27570 27806 27582 27858
rect 27634 27806 27646 27858
rect 26686 27794 26738 27806
rect 30046 27794 30098 27806
rect 2494 27746 2546 27758
rect 2494 27682 2546 27694
rect 3390 27746 3442 27758
rect 5406 27746 5458 27758
rect 22654 27746 22706 27758
rect 3938 27694 3950 27746
rect 4002 27694 4014 27746
rect 9986 27694 9998 27746
rect 10050 27694 10062 27746
rect 3390 27682 3442 27694
rect 5406 27682 5458 27694
rect 22654 27682 22706 27694
rect 24670 27746 24722 27758
rect 24670 27682 24722 27694
rect 28142 27746 28194 27758
rect 28142 27682 28194 27694
rect 29150 27746 29202 27758
rect 29150 27682 29202 27694
rect 16718 27634 16770 27646
rect 16258 27582 16270 27634
rect 16322 27582 16334 27634
rect 19282 27582 19294 27634
rect 19346 27582 19358 27634
rect 16718 27570 16770 27582
rect 1344 27466 58576 27500
rect 1344 27414 4478 27466
rect 4530 27414 4582 27466
rect 4634 27414 4686 27466
rect 4738 27414 35198 27466
rect 35250 27414 35302 27466
rect 35354 27414 35406 27466
rect 35458 27414 58576 27466
rect 1344 27380 58576 27414
rect 15822 27298 15874 27310
rect 24770 27246 24782 27298
rect 24834 27246 24846 27298
rect 15822 27234 15874 27246
rect 6414 27186 6466 27198
rect 6414 27122 6466 27134
rect 8878 27186 8930 27198
rect 8878 27122 8930 27134
rect 9214 27186 9266 27198
rect 9214 27122 9266 27134
rect 10558 27186 10610 27198
rect 10558 27122 10610 27134
rect 12686 27186 12738 27198
rect 12686 27122 12738 27134
rect 14142 27186 14194 27198
rect 14142 27122 14194 27134
rect 14478 27186 14530 27198
rect 14478 27122 14530 27134
rect 17166 27186 17218 27198
rect 17166 27122 17218 27134
rect 17502 27186 17554 27198
rect 17502 27122 17554 27134
rect 17950 27186 18002 27198
rect 17950 27122 18002 27134
rect 18398 27186 18450 27198
rect 18398 27122 18450 27134
rect 19294 27186 19346 27198
rect 19294 27122 19346 27134
rect 20190 27186 20242 27198
rect 20190 27122 20242 27134
rect 23774 27186 23826 27198
rect 23774 27122 23826 27134
rect 26574 27186 26626 27198
rect 26574 27122 26626 27134
rect 27134 27186 27186 27198
rect 27134 27122 27186 27134
rect 9102 27074 9154 27086
rect 5954 27022 5966 27074
rect 6018 27022 6030 27074
rect 9102 27010 9154 27022
rect 9774 27074 9826 27086
rect 13582 27074 13634 27086
rect 12226 27022 12238 27074
rect 12290 27022 12302 27074
rect 9774 27010 9826 27022
rect 13582 27010 13634 27022
rect 14702 27074 14754 27086
rect 14702 27010 14754 27022
rect 15374 27074 15426 27086
rect 15374 27010 15426 27022
rect 15710 27074 15762 27086
rect 15710 27010 15762 27022
rect 18510 27074 18562 27086
rect 26126 27074 26178 27086
rect 18834 27022 18846 27074
rect 18898 27022 18910 27074
rect 24210 27022 24222 27074
rect 24274 27022 24286 27074
rect 24434 27022 24446 27074
rect 24498 27022 24510 27074
rect 25218 27022 25230 27074
rect 25282 27022 25294 27074
rect 18510 27010 18562 27022
rect 26126 27010 26178 27022
rect 4734 26962 4786 26974
rect 4734 26898 4786 26910
rect 10110 26962 10162 26974
rect 10110 26898 10162 26910
rect 15150 26962 15202 26974
rect 15150 26898 15202 26910
rect 15262 26962 15314 26974
rect 15262 26898 15314 26910
rect 18286 26962 18338 26974
rect 25778 26910 25790 26962
rect 25842 26910 25854 26962
rect 18286 26898 18338 26910
rect 9326 26850 9378 26862
rect 9326 26786 9378 26798
rect 15822 26850 15874 26862
rect 15822 26786 15874 26798
rect 16606 26850 16658 26862
rect 16606 26786 16658 26798
rect 21870 26850 21922 26862
rect 21870 26786 21922 26798
rect 1344 26682 58576 26716
rect 1344 26630 19838 26682
rect 19890 26630 19942 26682
rect 19994 26630 20046 26682
rect 20098 26630 50558 26682
rect 50610 26630 50662 26682
rect 50714 26630 50766 26682
rect 50818 26630 58576 26682
rect 1344 26596 58576 26630
rect 6974 26514 7026 26526
rect 6974 26450 7026 26462
rect 7310 26514 7362 26526
rect 7310 26450 7362 26462
rect 9662 26514 9714 26526
rect 9662 26450 9714 26462
rect 9774 26514 9826 26526
rect 9774 26450 9826 26462
rect 10558 26514 10610 26526
rect 10558 26450 10610 26462
rect 12798 26514 12850 26526
rect 12798 26450 12850 26462
rect 13246 26514 13298 26526
rect 13246 26450 13298 26462
rect 13694 26514 13746 26526
rect 13694 26450 13746 26462
rect 14702 26514 14754 26526
rect 14702 26450 14754 26462
rect 15038 26514 15090 26526
rect 15038 26450 15090 26462
rect 15598 26514 15650 26526
rect 15598 26450 15650 26462
rect 15710 26514 15762 26526
rect 15710 26450 15762 26462
rect 17726 26514 17778 26526
rect 17726 26450 17778 26462
rect 25902 26514 25954 26526
rect 25902 26450 25954 26462
rect 26462 26514 26514 26526
rect 26462 26450 26514 26462
rect 7870 26402 7922 26414
rect 7870 26338 7922 26350
rect 11006 26402 11058 26414
rect 11006 26338 11058 26350
rect 15374 26402 15426 26414
rect 15374 26338 15426 26350
rect 17614 26402 17666 26414
rect 17614 26338 17666 26350
rect 18510 26402 18562 26414
rect 18510 26338 18562 26350
rect 5518 26290 5570 26302
rect 9550 26290 9602 26302
rect 5954 26238 5966 26290
rect 6018 26238 6030 26290
rect 5518 26226 5570 26238
rect 9550 26226 9602 26238
rect 10222 26290 10274 26302
rect 10222 26226 10274 26238
rect 11342 26290 11394 26302
rect 11342 26226 11394 26238
rect 11902 26290 11954 26302
rect 11902 26226 11954 26238
rect 12238 26290 12290 26302
rect 12238 26226 12290 26238
rect 15822 26290 15874 26302
rect 17838 26290 17890 26302
rect 16034 26238 16046 26290
rect 16098 26238 16110 26290
rect 17378 26238 17390 26290
rect 17442 26238 17454 26290
rect 15822 26226 15874 26238
rect 17838 26226 17890 26238
rect 17950 26290 18002 26302
rect 17950 26226 18002 26238
rect 21086 26290 21138 26302
rect 21086 26226 21138 26238
rect 21646 26290 21698 26302
rect 21646 26226 21698 26238
rect 22094 26290 22146 26302
rect 22094 26226 22146 26238
rect 14142 26178 14194 26190
rect 14142 26114 14194 26126
rect 16830 26178 16882 26190
rect 16830 26114 16882 26126
rect 19070 26178 19122 26190
rect 19070 26114 19122 26126
rect 19854 26178 19906 26190
rect 19854 26114 19906 26126
rect 20302 26178 20354 26190
rect 20302 26114 20354 26126
rect 20750 26178 20802 26190
rect 20750 26114 20802 26126
rect 22654 26178 22706 26190
rect 22654 26114 22706 26126
rect 23102 26178 23154 26190
rect 25442 26126 25454 26178
rect 25506 26126 25518 26178
rect 23102 26114 23154 26126
rect 1344 25898 58576 25932
rect 1344 25846 4478 25898
rect 4530 25846 4582 25898
rect 4634 25846 4686 25898
rect 4738 25846 35198 25898
rect 35250 25846 35302 25898
rect 35354 25846 35406 25898
rect 35458 25846 58576 25898
rect 1344 25812 58576 25846
rect 7310 25730 7362 25742
rect 7310 25666 7362 25678
rect 7086 25618 7138 25630
rect 23438 25618 23490 25630
rect 8642 25566 8654 25618
rect 8706 25566 8718 25618
rect 13906 25566 13918 25618
rect 13970 25566 13982 25618
rect 16482 25566 16494 25618
rect 16546 25566 16558 25618
rect 17714 25566 17726 25618
rect 17778 25566 17790 25618
rect 18050 25566 18062 25618
rect 18114 25566 18126 25618
rect 19954 25566 19966 25618
rect 20018 25566 20030 25618
rect 7086 25554 7138 25566
rect 23438 25554 23490 25566
rect 27134 25618 27186 25630
rect 28242 25566 28254 25618
rect 28306 25566 28318 25618
rect 27134 25554 27186 25566
rect 7534 25506 7586 25518
rect 7534 25442 7586 25454
rect 7646 25506 7698 25518
rect 9438 25506 9490 25518
rect 8978 25454 8990 25506
rect 9042 25454 9054 25506
rect 7646 25442 7698 25454
rect 9438 25442 9490 25454
rect 9662 25506 9714 25518
rect 9662 25442 9714 25454
rect 10222 25506 10274 25518
rect 10222 25442 10274 25454
rect 10446 25506 10498 25518
rect 11790 25506 11842 25518
rect 10994 25454 11006 25506
rect 11058 25454 11070 25506
rect 10446 25442 10498 25454
rect 11790 25442 11842 25454
rect 11902 25506 11954 25518
rect 11902 25442 11954 25454
rect 12014 25506 12066 25518
rect 12910 25506 12962 25518
rect 12338 25454 12350 25506
rect 12402 25454 12414 25506
rect 14466 25454 14478 25506
rect 14530 25454 14542 25506
rect 15586 25454 15598 25506
rect 15650 25454 15662 25506
rect 16034 25454 16046 25506
rect 16098 25454 16110 25506
rect 17378 25454 17390 25506
rect 17442 25454 17454 25506
rect 18386 25454 18398 25506
rect 18450 25454 18462 25506
rect 18834 25454 18846 25506
rect 18898 25454 18910 25506
rect 19730 25454 19742 25506
rect 19794 25454 19806 25506
rect 20066 25454 20078 25506
rect 20130 25454 20142 25506
rect 21746 25454 21758 25506
rect 21810 25454 21822 25506
rect 23650 25454 23662 25506
rect 23714 25454 23726 25506
rect 25330 25454 25342 25506
rect 25394 25454 25406 25506
rect 25554 25454 25566 25506
rect 25618 25454 25630 25506
rect 12014 25442 12066 25454
rect 12910 25442 12962 25454
rect 1710 25394 1762 25406
rect 1710 25330 1762 25342
rect 2046 25394 2098 25406
rect 2046 25330 2098 25342
rect 2494 25394 2546 25406
rect 2494 25330 2546 25342
rect 7870 25394 7922 25406
rect 7870 25330 7922 25342
rect 9550 25394 9602 25406
rect 9550 25330 9602 25342
rect 10782 25394 10834 25406
rect 10782 25330 10834 25342
rect 12574 25394 12626 25406
rect 14690 25342 14702 25394
rect 14754 25342 14766 25394
rect 16258 25342 16270 25394
rect 16322 25342 16334 25394
rect 20402 25342 20414 25394
rect 20466 25342 20478 25394
rect 22418 25342 22430 25394
rect 22482 25342 22494 25394
rect 23538 25342 23550 25394
rect 23602 25342 23614 25394
rect 12574 25330 12626 25342
rect 9886 25282 9938 25294
rect 12798 25282 12850 25294
rect 11330 25230 11342 25282
rect 11394 25230 11406 25282
rect 9886 25218 9938 25230
rect 12798 25218 12850 25230
rect 13470 25282 13522 25294
rect 21534 25282 21586 25294
rect 15250 25230 15262 25282
rect 15314 25230 15326 25282
rect 18610 25230 18622 25282
rect 18674 25230 18686 25282
rect 13470 25218 13522 25230
rect 21534 25218 21586 25230
rect 27806 25282 27858 25294
rect 27806 25218 27858 25230
rect 29262 25282 29314 25294
rect 29262 25218 29314 25230
rect 1344 25114 58576 25148
rect 1344 25062 19838 25114
rect 19890 25062 19942 25114
rect 19994 25062 20046 25114
rect 20098 25062 50558 25114
rect 50610 25062 50662 25114
rect 50714 25062 50766 25114
rect 50818 25062 58576 25114
rect 1344 25028 58576 25062
rect 6974 24946 7026 24958
rect 6974 24882 7026 24894
rect 7198 24946 7250 24958
rect 7198 24882 7250 24894
rect 8318 24946 8370 24958
rect 8318 24882 8370 24894
rect 11230 24946 11282 24958
rect 11230 24882 11282 24894
rect 11678 24946 11730 24958
rect 17614 24946 17666 24958
rect 25790 24946 25842 24958
rect 16706 24894 16718 24946
rect 16770 24894 16782 24946
rect 22754 24894 22766 24946
rect 22818 24894 22830 24946
rect 11678 24882 11730 24894
rect 17614 24882 17666 24894
rect 25790 24882 25842 24894
rect 26238 24946 26290 24958
rect 26238 24882 26290 24894
rect 16034 24782 16046 24834
rect 16098 24782 16110 24834
rect 19282 24782 19294 24834
rect 19346 24782 19358 24834
rect 20402 24782 20414 24834
rect 20466 24782 20478 24834
rect 22082 24782 22094 24834
rect 22146 24782 22158 24834
rect 24210 24782 24222 24834
rect 24274 24782 24286 24834
rect 7758 24722 7810 24734
rect 12898 24670 12910 24722
rect 12962 24670 12974 24722
rect 13346 24670 13358 24722
rect 13410 24670 13422 24722
rect 13570 24670 13582 24722
rect 13634 24670 13646 24722
rect 13906 24670 13918 24722
rect 13970 24670 13982 24722
rect 16482 24670 16494 24722
rect 16546 24670 16558 24722
rect 17826 24670 17838 24722
rect 17890 24670 17902 24722
rect 21074 24670 21086 24722
rect 21138 24670 21150 24722
rect 22306 24670 22318 24722
rect 22370 24670 22382 24722
rect 24434 24670 24446 24722
rect 24498 24670 24510 24722
rect 7758 24658 7810 24670
rect 25230 24610 25282 24622
rect 18498 24558 18510 24610
rect 18562 24558 18574 24610
rect 25230 24546 25282 24558
rect 1344 24330 58576 24364
rect 1344 24278 4478 24330
rect 4530 24278 4582 24330
rect 4634 24278 4686 24330
rect 4738 24278 35198 24330
rect 35250 24278 35302 24330
rect 35354 24278 35406 24330
rect 35458 24278 58576 24330
rect 1344 24244 58576 24278
rect 20738 24110 20750 24162
rect 20802 24110 20814 24162
rect 11678 24050 11730 24062
rect 11678 23986 11730 23998
rect 13022 24050 13074 24062
rect 16158 24050 16210 24062
rect 23326 24050 23378 24062
rect 25230 24050 25282 24062
rect 14018 23998 14030 24050
rect 14082 23998 14094 24050
rect 15138 23998 15150 24050
rect 15202 23998 15214 24050
rect 19730 23998 19742 24050
rect 19794 23998 19806 24050
rect 21858 23998 21870 24050
rect 21922 23998 21934 24050
rect 24322 23998 24334 24050
rect 24386 23998 24398 24050
rect 13022 23986 13074 23998
rect 16158 23986 16210 23998
rect 23326 23986 23378 23998
rect 25230 23986 25282 23998
rect 25790 24050 25842 24062
rect 25790 23986 25842 23998
rect 20190 23938 20242 23950
rect 14690 23886 14702 23938
rect 14754 23886 14766 23938
rect 15474 23886 15486 23938
rect 15538 23886 15550 23938
rect 16370 23886 16382 23938
rect 16434 23886 16446 23938
rect 18050 23886 18062 23938
rect 18114 23886 18126 23938
rect 19954 23886 19966 23938
rect 20018 23886 20030 23938
rect 20190 23874 20242 23886
rect 20302 23938 20354 23950
rect 24782 23938 24834 23950
rect 21970 23886 21982 23938
rect 22034 23886 22046 23938
rect 22306 23886 22318 23938
rect 22370 23886 22382 23938
rect 23762 23886 23774 23938
rect 23826 23886 23838 23938
rect 20302 23874 20354 23886
rect 24782 23874 24834 23886
rect 1710 23826 1762 23838
rect 1710 23762 1762 23774
rect 2046 23826 2098 23838
rect 16930 23774 16942 23826
rect 16994 23774 17006 23826
rect 18162 23774 18174 23826
rect 18226 23774 18238 23826
rect 21298 23774 21310 23826
rect 21362 23774 21374 23826
rect 2046 23762 2098 23774
rect 2494 23714 2546 23726
rect 2494 23650 2546 23662
rect 1344 23546 58576 23580
rect 1344 23494 19838 23546
rect 19890 23494 19942 23546
rect 19994 23494 20046 23546
rect 20098 23494 50558 23546
rect 50610 23494 50662 23546
rect 50714 23494 50766 23546
rect 50818 23494 58576 23546
rect 1344 23460 58576 23494
rect 15598 23378 15650 23390
rect 15598 23314 15650 23326
rect 15934 23378 15986 23390
rect 15934 23314 15986 23326
rect 16158 23378 16210 23390
rect 16158 23314 16210 23326
rect 16718 23378 16770 23390
rect 16718 23314 16770 23326
rect 18622 23378 18674 23390
rect 18622 23314 18674 23326
rect 19070 23378 19122 23390
rect 19070 23314 19122 23326
rect 21086 23378 21138 23390
rect 21086 23314 21138 23326
rect 21646 23378 21698 23390
rect 21646 23314 21698 23326
rect 22206 23378 22258 23390
rect 22206 23314 22258 23326
rect 22990 23378 23042 23390
rect 22990 23314 23042 23326
rect 25454 23378 25506 23390
rect 25454 23314 25506 23326
rect 15822 23266 15874 23278
rect 15822 23202 15874 23214
rect 19182 23266 19234 23278
rect 21298 23214 21310 23266
rect 21362 23214 21374 23266
rect 19182 23202 19234 23214
rect 15150 23042 15202 23054
rect 15150 22978 15202 22990
rect 17614 23042 17666 23054
rect 17614 22978 17666 22990
rect 19070 22930 19122 22942
rect 19070 22866 19122 22878
rect 1344 22762 58576 22796
rect 1344 22710 4478 22762
rect 4530 22710 4582 22762
rect 4634 22710 4686 22762
rect 4738 22710 35198 22762
rect 35250 22710 35302 22762
rect 35354 22710 35406 22762
rect 35458 22710 58576 22762
rect 1344 22676 58576 22710
rect 15598 22482 15650 22494
rect 15598 22418 15650 22430
rect 1710 22258 1762 22270
rect 1710 22194 1762 22206
rect 2046 22258 2098 22270
rect 2046 22194 2098 22206
rect 2494 22146 2546 22158
rect 2494 22082 2546 22094
rect 1344 21978 58576 22012
rect 1344 21926 19838 21978
rect 19890 21926 19942 21978
rect 19994 21926 20046 21978
rect 20098 21926 50558 21978
rect 50610 21926 50662 21978
rect 50714 21926 50766 21978
rect 50818 21926 58576 21978
rect 1344 21892 58576 21926
rect 1344 21194 58576 21228
rect 1344 21142 4478 21194
rect 4530 21142 4582 21194
rect 4634 21142 4686 21194
rect 4738 21142 35198 21194
rect 35250 21142 35302 21194
rect 35354 21142 35406 21194
rect 35458 21142 58576 21194
rect 1344 21108 58576 21142
rect 2034 20638 2046 20690
rect 2098 20638 2110 20690
rect 1710 20578 1762 20590
rect 1710 20514 1762 20526
rect 2494 20578 2546 20590
rect 2494 20514 2546 20526
rect 1344 20410 58576 20444
rect 1344 20358 19838 20410
rect 19890 20358 19942 20410
rect 19994 20358 20046 20410
rect 20098 20358 50558 20410
rect 50610 20358 50662 20410
rect 50714 20358 50766 20410
rect 50818 20358 58576 20410
rect 1344 20324 58576 20358
rect 1344 19626 58576 19660
rect 1344 19574 4478 19626
rect 4530 19574 4582 19626
rect 4634 19574 4686 19626
rect 4738 19574 35198 19626
rect 35250 19574 35302 19626
rect 35354 19574 35406 19626
rect 35458 19574 58576 19626
rect 1344 19540 58576 19574
rect 1344 18842 58576 18876
rect 1344 18790 19838 18842
rect 19890 18790 19942 18842
rect 19994 18790 20046 18842
rect 20098 18790 50558 18842
rect 50610 18790 50662 18842
rect 50714 18790 50766 18842
rect 50818 18790 58576 18842
rect 1344 18756 58576 18790
rect 2046 18674 2098 18686
rect 2046 18610 2098 18622
rect 1710 18450 1762 18462
rect 1710 18386 1762 18398
rect 2494 18338 2546 18350
rect 2494 18274 2546 18286
rect 1344 18058 58576 18092
rect 1344 18006 4478 18058
rect 4530 18006 4582 18058
rect 4634 18006 4686 18058
rect 4738 18006 35198 18058
rect 35250 18006 35302 18058
rect 35354 18006 35406 18058
rect 35458 18006 58576 18058
rect 1344 17972 58576 18006
rect 1344 17274 58576 17308
rect 1344 17222 19838 17274
rect 19890 17222 19942 17274
rect 19994 17222 20046 17274
rect 20098 17222 50558 17274
rect 50610 17222 50662 17274
rect 50714 17222 50766 17274
rect 50818 17222 58576 17274
rect 1344 17188 58576 17222
rect 2034 17054 2046 17106
rect 2098 17054 2110 17106
rect 1710 16882 1762 16894
rect 1710 16818 1762 16830
rect 2494 16882 2546 16894
rect 2494 16818 2546 16830
rect 1344 16490 58576 16524
rect 1344 16438 4478 16490
rect 4530 16438 4582 16490
rect 4634 16438 4686 16490
rect 4738 16438 35198 16490
rect 35250 16438 35302 16490
rect 35354 16438 35406 16490
rect 35458 16438 58576 16490
rect 1344 16404 58576 16438
rect 1344 15706 58576 15740
rect 1344 15654 19838 15706
rect 19890 15654 19942 15706
rect 19994 15654 20046 15706
rect 20098 15654 50558 15706
rect 50610 15654 50662 15706
rect 50714 15654 50766 15706
rect 50818 15654 58576 15706
rect 1344 15620 58576 15654
rect 2046 15538 2098 15550
rect 2046 15474 2098 15486
rect 1710 15314 1762 15326
rect 1710 15250 1762 15262
rect 2494 15202 2546 15214
rect 2494 15138 2546 15150
rect 1344 14922 58576 14956
rect 1344 14870 4478 14922
rect 4530 14870 4582 14922
rect 4634 14870 4686 14922
rect 4738 14870 35198 14922
rect 35250 14870 35302 14922
rect 35354 14870 35406 14922
rect 35458 14870 58576 14922
rect 1344 14836 58576 14870
rect 1344 14138 58576 14172
rect 1344 14086 19838 14138
rect 19890 14086 19942 14138
rect 19994 14086 20046 14138
rect 20098 14086 50558 14138
rect 50610 14086 50662 14138
rect 50714 14086 50766 14138
rect 50818 14086 58576 14138
rect 1344 14052 58576 14086
rect 1344 13354 58576 13388
rect 1344 13302 4478 13354
rect 4530 13302 4582 13354
rect 4634 13302 4686 13354
rect 4738 13302 35198 13354
rect 35250 13302 35302 13354
rect 35354 13302 35406 13354
rect 35458 13302 58576 13354
rect 1344 13268 58576 13302
rect 1710 12850 1762 12862
rect 1710 12786 1762 12798
rect 2046 12850 2098 12862
rect 2046 12786 2098 12798
rect 2494 12850 2546 12862
rect 2494 12786 2546 12798
rect 1344 12570 58576 12604
rect 1344 12518 19838 12570
rect 19890 12518 19942 12570
rect 19994 12518 20046 12570
rect 20098 12518 50558 12570
rect 50610 12518 50662 12570
rect 50714 12518 50766 12570
rect 50818 12518 58576 12570
rect 1344 12484 58576 12518
rect 1344 11786 58576 11820
rect 1344 11734 4478 11786
rect 4530 11734 4582 11786
rect 4634 11734 4686 11786
rect 4738 11734 35198 11786
rect 35250 11734 35302 11786
rect 35354 11734 35406 11786
rect 35458 11734 58576 11786
rect 1344 11700 58576 11734
rect 1710 11282 1762 11294
rect 1710 11218 1762 11230
rect 2046 11282 2098 11294
rect 2046 11218 2098 11230
rect 2494 11170 2546 11182
rect 2494 11106 2546 11118
rect 1344 11002 58576 11036
rect 1344 10950 19838 11002
rect 19890 10950 19942 11002
rect 19994 10950 20046 11002
rect 20098 10950 50558 11002
rect 50610 10950 50662 11002
rect 50714 10950 50766 11002
rect 50818 10950 58576 11002
rect 1344 10916 58576 10950
rect 1344 10218 58576 10252
rect 1344 10166 4478 10218
rect 4530 10166 4582 10218
rect 4634 10166 4686 10218
rect 4738 10166 35198 10218
rect 35250 10166 35302 10218
rect 35354 10166 35406 10218
rect 35458 10166 58576 10218
rect 1344 10132 58576 10166
rect 1710 9714 1762 9726
rect 1710 9650 1762 9662
rect 2046 9714 2098 9726
rect 2046 9650 2098 9662
rect 2494 9602 2546 9614
rect 2494 9538 2546 9550
rect 1344 9434 58576 9468
rect 1344 9382 19838 9434
rect 19890 9382 19942 9434
rect 19994 9382 20046 9434
rect 20098 9382 50558 9434
rect 50610 9382 50662 9434
rect 50714 9382 50766 9434
rect 50818 9382 58576 9434
rect 1344 9348 58576 9382
rect 1344 8650 58576 8684
rect 1344 8598 4478 8650
rect 4530 8598 4582 8650
rect 4634 8598 4686 8650
rect 4738 8598 35198 8650
rect 35250 8598 35302 8650
rect 35354 8598 35406 8650
rect 35458 8598 58576 8650
rect 1344 8564 58576 8598
rect 1710 8146 1762 8158
rect 1710 8082 1762 8094
rect 2046 8146 2098 8158
rect 2046 8082 2098 8094
rect 2494 8034 2546 8046
rect 2494 7970 2546 7982
rect 1344 7866 58576 7900
rect 1344 7814 19838 7866
rect 19890 7814 19942 7866
rect 19994 7814 20046 7866
rect 20098 7814 50558 7866
rect 50610 7814 50662 7866
rect 50714 7814 50766 7866
rect 50818 7814 58576 7866
rect 1344 7780 58576 7814
rect 1344 7082 58576 7116
rect 1344 7030 4478 7082
rect 4530 7030 4582 7082
rect 4634 7030 4686 7082
rect 4738 7030 35198 7082
rect 35250 7030 35302 7082
rect 35354 7030 35406 7082
rect 35458 7030 58576 7082
rect 1344 6996 58576 7030
rect 1344 6298 58576 6332
rect 1344 6246 19838 6298
rect 19890 6246 19942 6298
rect 19994 6246 20046 6298
rect 20098 6246 50558 6298
rect 50610 6246 50662 6298
rect 50714 6246 50766 6298
rect 50818 6246 58576 6298
rect 1344 6212 58576 6246
rect 1710 5906 1762 5918
rect 1710 5842 1762 5854
rect 2146 5742 2158 5794
rect 2210 5742 2222 5794
rect 1344 5514 58576 5548
rect 1344 5462 4478 5514
rect 4530 5462 4582 5514
rect 4634 5462 4686 5514
rect 4738 5462 35198 5514
rect 35250 5462 35302 5514
rect 35354 5462 35406 5514
rect 35458 5462 58576 5514
rect 1344 5428 58576 5462
rect 1822 5234 1874 5246
rect 1822 5170 1874 5182
rect 1344 4730 58576 4764
rect 1344 4678 19838 4730
rect 19890 4678 19942 4730
rect 19994 4678 20046 4730
rect 20098 4678 50558 4730
rect 50610 4678 50662 4730
rect 50714 4678 50766 4730
rect 50818 4678 58576 4730
rect 1344 4644 58576 4678
rect 2046 4562 2098 4574
rect 2046 4498 2098 4510
rect 1710 4338 1762 4350
rect 1710 4274 1762 4286
rect 2494 4226 2546 4238
rect 2494 4162 2546 4174
rect 1344 3946 58576 3980
rect 1344 3894 4478 3946
rect 4530 3894 4582 3946
rect 4634 3894 4686 3946
rect 4738 3894 35198 3946
rect 35250 3894 35302 3946
rect 35354 3894 35406 3946
rect 35458 3894 58576 3946
rect 1344 3860 58576 3894
rect 2270 3666 2322 3678
rect 2270 3602 2322 3614
rect 1710 3442 1762 3454
rect 1710 3378 1762 3390
rect 2718 3442 2770 3454
rect 2718 3378 2770 3390
rect 1344 3162 58576 3196
rect 1344 3110 19838 3162
rect 19890 3110 19942 3162
rect 19994 3110 20046 3162
rect 20098 3110 50558 3162
rect 50610 3110 50662 3162
rect 50714 3110 50766 3162
rect 50818 3110 58576 3162
rect 1344 3076 58576 3110
<< via1 >>
rect 38782 56590 38834 56642
rect 39342 56590 39394 56642
rect 40126 56590 40178 56642
rect 19838 56422 19890 56474
rect 19942 56422 19994 56474
rect 20046 56422 20098 56474
rect 50558 56422 50610 56474
rect 50662 56422 50714 56474
rect 50766 56422 50818 56474
rect 5070 56254 5122 56306
rect 7422 56254 7474 56306
rect 7646 56254 7698 56306
rect 9662 56254 9714 56306
rect 9886 56254 9938 56306
rect 11902 56254 11954 56306
rect 12126 56254 12178 56306
rect 14142 56254 14194 56306
rect 16494 56254 16546 56306
rect 16942 56254 16994 56306
rect 18622 56254 18674 56306
rect 18846 56254 18898 56306
rect 20302 56254 20354 56306
rect 23102 56254 23154 56306
rect 25342 56254 25394 56306
rect 27918 56254 27970 56306
rect 29822 56254 29874 56306
rect 31726 56254 31778 56306
rect 34302 56254 34354 56306
rect 36542 56254 36594 56306
rect 39342 56254 39394 56306
rect 41470 56254 41522 56306
rect 44606 56254 44658 56306
rect 48974 56254 49026 56306
rect 52222 56254 52274 56306
rect 56030 56254 56082 56306
rect 2046 56142 2098 56194
rect 2382 56142 2434 56194
rect 5518 56142 5570 56194
rect 5854 56142 5906 56194
rect 7982 56142 8034 56194
rect 10222 56142 10274 56194
rect 12462 56142 12514 56194
rect 14366 56142 14418 56194
rect 17278 56142 17330 56194
rect 19182 56142 19234 56194
rect 21086 56142 21138 56194
rect 21422 56142 21474 56194
rect 23326 56142 23378 56194
rect 25566 56142 25618 56194
rect 28366 56142 28418 56194
rect 30046 56142 30098 56194
rect 32286 56142 32338 56194
rect 32622 56142 32674 56194
rect 34526 56142 34578 56194
rect 34862 56142 34914 56194
rect 36766 56142 36818 56194
rect 37102 56142 37154 56194
rect 39790 56142 39842 56194
rect 40126 56142 40178 56194
rect 1710 56030 1762 56082
rect 2606 56030 2658 56082
rect 14590 56030 14642 56082
rect 23550 56030 23602 56082
rect 25790 56030 25842 56082
rect 28590 56030 28642 56082
rect 30270 56030 30322 56082
rect 40462 56030 40514 56082
rect 43710 56030 43762 56082
rect 47742 56030 47794 56082
rect 47966 56030 48018 56082
rect 51214 56030 51266 56082
rect 54574 56030 54626 56082
rect 55022 56030 55074 56082
rect 3166 55918 3218 55970
rect 37998 55918 38050 55970
rect 38894 55918 38946 55970
rect 4478 55638 4530 55690
rect 4582 55638 4634 55690
rect 4686 55638 4738 55690
rect 35198 55638 35250 55690
rect 35302 55638 35354 55690
rect 35406 55638 35458 55690
rect 2158 55358 2210 55410
rect 16382 55358 16434 55410
rect 20526 55358 20578 55410
rect 32062 55358 32114 55410
rect 36430 55358 36482 55410
rect 39230 55358 39282 55410
rect 43150 55358 43202 55410
rect 46734 55358 46786 55410
rect 53678 55358 53730 55410
rect 56702 55358 56754 55410
rect 13582 55246 13634 55298
rect 16830 55246 16882 55298
rect 17726 55246 17778 55298
rect 21422 55246 21474 55298
rect 22990 55246 23042 55298
rect 25342 55246 25394 55298
rect 27694 55246 27746 55298
rect 29262 55246 29314 55298
rect 32622 55246 32674 55298
rect 33182 55246 33234 55298
rect 33630 55246 33682 55298
rect 37102 55246 37154 55298
rect 40350 55246 40402 55298
rect 45726 55246 45778 55298
rect 52670 55246 52722 55298
rect 55582 55246 55634 55298
rect 11790 55134 11842 55186
rect 14254 55134 14306 55186
rect 18398 55134 18450 55186
rect 29934 55134 29986 55186
rect 34302 55134 34354 55186
rect 37326 55134 37378 55186
rect 41022 55134 41074 55186
rect 11902 55022 11954 55074
rect 22878 55022 22930 55074
rect 25230 55022 25282 55074
rect 27582 55022 27634 55074
rect 32622 55022 32674 55074
rect 37774 55022 37826 55074
rect 38222 55022 38274 55074
rect 38558 55022 38610 55074
rect 39118 55022 39170 55074
rect 39902 55022 39954 55074
rect 43598 55022 43650 55074
rect 45390 55022 45442 55074
rect 50878 55022 50930 55074
rect 52110 55022 52162 55074
rect 19838 54854 19890 54906
rect 19942 54854 19994 54906
rect 20046 54854 20098 54906
rect 50558 54854 50610 54906
rect 50662 54854 50714 54906
rect 50766 54854 50818 54906
rect 12462 54686 12514 54738
rect 14814 54686 14866 54738
rect 15822 54686 15874 54738
rect 17614 54686 17666 54738
rect 18510 54686 18562 54738
rect 29934 54686 29986 54738
rect 33966 54686 34018 54738
rect 36430 54686 36482 54738
rect 40350 54686 40402 54738
rect 40910 54686 40962 54738
rect 2046 54574 2098 54626
rect 12798 54574 12850 54626
rect 13246 54574 13298 54626
rect 15262 54574 15314 54626
rect 18734 54574 18786 54626
rect 29150 54574 29202 54626
rect 29486 54574 29538 54626
rect 31838 54574 31890 54626
rect 34750 54574 34802 54626
rect 36654 54574 36706 54626
rect 38894 54574 38946 54626
rect 41694 54574 41746 54626
rect 1710 54462 1762 54514
rect 13694 54462 13746 54514
rect 14590 54462 14642 54514
rect 15038 54462 15090 54514
rect 15710 54462 15762 54514
rect 15934 54462 15986 54514
rect 16382 54462 16434 54514
rect 17278 54462 17330 54514
rect 17726 54462 17778 54514
rect 17838 54462 17890 54514
rect 18286 54462 18338 54514
rect 18398 54462 18450 54514
rect 21086 54462 21138 54514
rect 25342 54462 25394 54514
rect 28814 54462 28866 54514
rect 29822 54462 29874 54514
rect 30046 54462 30098 54514
rect 30606 54462 30658 54514
rect 33182 54462 33234 54514
rect 33406 54462 33458 54514
rect 33966 54462 34018 54514
rect 38558 54462 38610 54514
rect 41022 54462 41074 54514
rect 41358 54462 41410 54514
rect 2494 54350 2546 54402
rect 13806 54350 13858 54402
rect 21758 54350 21810 54402
rect 23886 54350 23938 54402
rect 26014 54350 26066 54402
rect 28142 54350 28194 54402
rect 31726 54350 31778 54402
rect 32510 54350 32562 54402
rect 34414 54350 34466 54402
rect 36318 54350 36370 54402
rect 38222 54350 38274 54402
rect 55246 54350 55298 54402
rect 30382 54238 30434 54290
rect 32062 54238 32114 54290
rect 33630 54238 33682 54290
rect 41246 54238 41298 54290
rect 4478 54070 4530 54122
rect 4582 54070 4634 54122
rect 4686 54070 4738 54122
rect 35198 54070 35250 54122
rect 35302 54070 35354 54122
rect 35406 54070 35458 54122
rect 40910 53902 40962 53954
rect 23662 53790 23714 53842
rect 29262 53790 29314 53842
rect 41022 53790 41074 53842
rect 42142 53790 42194 53842
rect 22430 53678 22482 53730
rect 22654 53678 22706 53730
rect 22878 53678 22930 53730
rect 23774 53678 23826 53730
rect 24558 53678 24610 53730
rect 33070 53678 33122 53730
rect 38334 53678 38386 53730
rect 41246 53678 41298 53730
rect 22318 53566 22370 53618
rect 25006 53566 25058 53618
rect 25230 53566 25282 53618
rect 26350 53566 26402 53618
rect 32622 53566 32674 53618
rect 33294 53566 33346 53618
rect 37774 53566 37826 53618
rect 38782 53566 38834 53618
rect 39118 53566 39170 53618
rect 42478 53566 42530 53618
rect 10446 53454 10498 53506
rect 11566 53454 11618 53506
rect 15486 53454 15538 53506
rect 16046 53454 16098 53506
rect 16382 53454 16434 53506
rect 16718 53454 16770 53506
rect 18174 53454 18226 53506
rect 21982 53454 22034 53506
rect 23550 53454 23602 53506
rect 23998 53454 24050 53506
rect 24894 53454 24946 53506
rect 25678 53454 25730 53506
rect 26238 53454 26290 53506
rect 26462 53454 26514 53506
rect 26686 53454 26738 53506
rect 38110 53454 38162 53506
rect 42254 53454 42306 53506
rect 19838 53286 19890 53338
rect 19942 53286 19994 53338
rect 20046 53286 20098 53338
rect 50558 53286 50610 53338
rect 50662 53286 50714 53338
rect 50766 53286 50818 53338
rect 12798 53118 12850 53170
rect 23438 53118 23490 53170
rect 29262 53118 29314 53170
rect 32062 53118 32114 53170
rect 33966 53118 34018 53170
rect 38446 53118 38498 53170
rect 41022 53118 41074 53170
rect 2046 53006 2098 53058
rect 9886 53006 9938 53058
rect 10558 53006 10610 53058
rect 12014 53006 12066 53058
rect 12350 53006 12402 53058
rect 22766 53006 22818 53058
rect 26686 53006 26738 53058
rect 29710 53006 29762 53058
rect 30046 53006 30098 53058
rect 30270 53006 30322 53058
rect 32286 53006 32338 53058
rect 36654 53006 36706 53058
rect 36766 53006 36818 53058
rect 1710 52894 1762 52946
rect 7982 52894 8034 52946
rect 8766 52894 8818 52946
rect 10222 52894 10274 52946
rect 10670 52894 10722 52946
rect 10894 52894 10946 52946
rect 11342 52894 11394 52946
rect 18062 52894 18114 52946
rect 18398 52894 18450 52946
rect 18510 52894 18562 52946
rect 22430 52894 22482 52946
rect 22990 52894 23042 52946
rect 25454 52894 25506 52946
rect 25902 52894 25954 52946
rect 26126 52894 26178 52946
rect 27022 52894 27074 52946
rect 30494 52894 30546 52946
rect 30830 52894 30882 52946
rect 33182 52894 33234 52946
rect 33406 52894 33458 52946
rect 33630 52894 33682 52946
rect 33966 52894 34018 52946
rect 36542 52894 36594 52946
rect 36990 52894 37042 52946
rect 37774 52894 37826 52946
rect 37998 52894 38050 52946
rect 41918 52894 41970 52946
rect 42702 52894 42754 52946
rect 2494 52782 2546 52834
rect 5854 52782 5906 52834
rect 15374 52782 15426 52834
rect 18174 52782 18226 52834
rect 19070 52782 19122 52834
rect 22542 52782 22594 52834
rect 26014 52782 26066 52834
rect 27470 52782 27522 52834
rect 30158 52782 30210 52834
rect 31950 52782 32002 52834
rect 37662 52782 37714 52834
rect 41582 52782 41634 52834
rect 44830 52782 44882 52834
rect 11006 52670 11058 52722
rect 29598 52670 29650 52722
rect 37438 52670 37490 52722
rect 41022 52670 41074 52722
rect 41470 52670 41522 52722
rect 4478 52502 4530 52554
rect 4582 52502 4634 52554
rect 4686 52502 4738 52554
rect 35198 52502 35250 52554
rect 35302 52502 35354 52554
rect 35406 52502 35458 52554
rect 10446 52334 10498 52386
rect 11678 52334 11730 52386
rect 12014 52334 12066 52386
rect 13022 52334 13074 52386
rect 41694 52334 41746 52386
rect 12798 52222 12850 52274
rect 17838 52222 17890 52274
rect 19966 52222 20018 52274
rect 30158 52222 30210 52274
rect 32286 52222 32338 52274
rect 32846 52222 32898 52274
rect 34190 52222 34242 52274
rect 36318 52222 36370 52274
rect 38670 52222 38722 52274
rect 42702 52222 42754 52274
rect 8990 52110 9042 52162
rect 9998 52110 10050 52162
rect 10334 52110 10386 52162
rect 10782 52110 10834 52162
rect 11118 52110 11170 52162
rect 11342 52110 11394 52162
rect 11902 52110 11954 52162
rect 12350 52110 12402 52162
rect 14590 52110 14642 52162
rect 14814 52110 14866 52162
rect 15598 52110 15650 52162
rect 16270 52110 16322 52162
rect 20638 52110 20690 52162
rect 27246 52110 27298 52162
rect 27694 52110 27746 52162
rect 29374 52110 29426 52162
rect 33518 52110 33570 52162
rect 38334 52110 38386 52162
rect 40238 52110 40290 52162
rect 41470 52110 41522 52162
rect 41918 52110 41970 52162
rect 42590 52110 42642 52162
rect 43038 52110 43090 52162
rect 15150 51998 15202 52050
rect 25230 51998 25282 52050
rect 39230 51998 39282 52050
rect 41246 51998 41298 52050
rect 41358 51998 41410 52050
rect 42254 51998 42306 52050
rect 10110 51886 10162 51938
rect 11902 51886 11954 51938
rect 14702 51886 14754 51938
rect 15710 51886 15762 51938
rect 15822 51886 15874 51938
rect 37102 51886 37154 51938
rect 19838 51718 19890 51770
rect 19942 51718 19994 51770
rect 20046 51718 20098 51770
rect 50558 51718 50610 51770
rect 50662 51718 50714 51770
rect 50766 51718 50818 51770
rect 12014 51550 12066 51602
rect 16494 51550 16546 51602
rect 17390 51550 17442 51602
rect 18174 51550 18226 51602
rect 18286 51550 18338 51602
rect 18622 51550 18674 51602
rect 40014 51550 40066 51602
rect 41806 51550 41858 51602
rect 42254 51550 42306 51602
rect 2046 51438 2098 51490
rect 10670 51438 10722 51490
rect 10894 51438 10946 51490
rect 13918 51438 13970 51490
rect 21758 51438 21810 51490
rect 40238 51438 40290 51490
rect 41022 51438 41074 51490
rect 41246 51438 41298 51490
rect 1822 51326 1874 51378
rect 4398 51326 4450 51378
rect 7646 51326 7698 51378
rect 11118 51326 11170 51378
rect 11230 51326 11282 51378
rect 13246 51326 13298 51378
rect 16830 51326 16882 51378
rect 17726 51326 17778 51378
rect 18398 51326 18450 51378
rect 21086 51326 21138 51378
rect 25342 51326 25394 51378
rect 38446 51326 38498 51378
rect 38782 51326 38834 51378
rect 39006 51326 39058 51378
rect 39566 51326 39618 51378
rect 41806 51326 41858 51378
rect 2494 51214 2546 51266
rect 5070 51214 5122 51266
rect 7198 51214 7250 51266
rect 10782 51214 10834 51266
rect 16046 51214 16098 51266
rect 23886 51214 23938 51266
rect 26126 51214 26178 51266
rect 28254 51214 28306 51266
rect 38894 51214 38946 51266
rect 39902 51214 39954 51266
rect 42142 51214 42194 51266
rect 39230 51102 39282 51154
rect 41582 51102 41634 51154
rect 42478 51102 42530 51154
rect 4478 50934 4530 50986
rect 4582 50934 4634 50986
rect 4686 50934 4738 50986
rect 35198 50934 35250 50986
rect 35302 50934 35354 50986
rect 35406 50934 35458 50986
rect 7310 50766 7362 50818
rect 1710 50654 1762 50706
rect 3838 50654 3890 50706
rect 5070 50654 5122 50706
rect 7086 50654 7138 50706
rect 15934 50654 15986 50706
rect 16494 50654 16546 50706
rect 23662 50654 23714 50706
rect 26462 50654 26514 50706
rect 27358 50654 27410 50706
rect 34526 50654 34578 50706
rect 37886 50654 37938 50706
rect 40014 50654 40066 50706
rect 40462 50654 40514 50706
rect 40910 50654 40962 50706
rect 42030 50654 42082 50706
rect 44158 50654 44210 50706
rect 4622 50542 4674 50594
rect 21870 50542 21922 50594
rect 22094 50542 22146 50594
rect 23774 50542 23826 50594
rect 24446 50542 24498 50594
rect 26238 50542 26290 50594
rect 26686 50542 26738 50594
rect 26798 50542 26850 50594
rect 30382 50542 30434 50594
rect 35086 50542 35138 50594
rect 37102 50542 37154 50594
rect 41246 50542 41298 50594
rect 18174 50430 18226 50482
rect 22430 50430 22482 50482
rect 23550 50430 23602 50482
rect 23998 50430 24050 50482
rect 24782 50430 24834 50482
rect 7646 50318 7698 50370
rect 11902 50318 11954 50370
rect 12574 50318 12626 50370
rect 16046 50318 16098 50370
rect 18286 50318 18338 50370
rect 18510 50318 18562 50370
rect 30718 50318 30770 50370
rect 32398 50318 32450 50370
rect 34862 50318 34914 50370
rect 19838 50150 19890 50202
rect 19942 50150 19994 50202
rect 20046 50150 20098 50202
rect 50558 50150 50610 50202
rect 50662 50150 50714 50202
rect 50766 50150 50818 50202
rect 5070 49982 5122 50034
rect 7086 49982 7138 50034
rect 11342 49982 11394 50034
rect 12014 49982 12066 50034
rect 13134 49982 13186 50034
rect 33070 49982 33122 50034
rect 41022 49982 41074 50034
rect 3838 49870 3890 49922
rect 7198 49870 7250 49922
rect 7534 49870 7586 49922
rect 17614 49870 17666 49922
rect 25230 49870 25282 49922
rect 27582 49870 27634 49922
rect 4622 49758 4674 49810
rect 6526 49758 6578 49810
rect 8430 49758 8482 49810
rect 8990 49758 9042 49810
rect 10558 49758 10610 49810
rect 11566 49758 11618 49810
rect 12238 49758 12290 49810
rect 12910 49758 12962 49810
rect 22654 49758 22706 49810
rect 23102 49758 23154 49810
rect 32174 49758 32226 49810
rect 33294 49758 33346 49810
rect 33742 49758 33794 49810
rect 34414 49758 34466 49810
rect 34750 49758 34802 49810
rect 35086 49758 35138 49810
rect 1710 49646 1762 49698
rect 8094 49646 8146 49698
rect 10110 49646 10162 49698
rect 24110 49646 24162 49698
rect 29262 49646 29314 49698
rect 31390 49646 31442 49698
rect 33182 49646 33234 49698
rect 34862 49646 34914 49698
rect 35422 49646 35474 49698
rect 6414 49534 6466 49586
rect 11230 49534 11282 49586
rect 11902 49534 11954 49586
rect 25342 49534 25394 49586
rect 27694 49534 27746 49586
rect 4478 49366 4530 49418
rect 4582 49366 4634 49418
rect 4686 49366 4738 49418
rect 35198 49366 35250 49418
rect 35302 49366 35354 49418
rect 35406 49366 35458 49418
rect 11118 49198 11170 49250
rect 15822 49198 15874 49250
rect 18734 49198 18786 49250
rect 10222 49086 10274 49138
rect 11342 49086 11394 49138
rect 11902 49086 11954 49138
rect 15486 49086 15538 49138
rect 19070 49086 19122 49138
rect 24558 49086 24610 49138
rect 29598 49086 29650 49138
rect 32958 49086 33010 49138
rect 33518 49086 33570 49138
rect 35646 49086 35698 49138
rect 6526 48974 6578 49026
rect 6974 48974 7026 49026
rect 11454 48974 11506 49026
rect 15374 48974 15426 49026
rect 18174 48974 18226 49026
rect 21870 48974 21922 49026
rect 22094 48974 22146 49026
rect 22206 48974 22258 49026
rect 24670 48974 24722 49026
rect 25566 48974 25618 49026
rect 27246 48974 27298 49026
rect 32510 48974 32562 49026
rect 36430 48974 36482 49026
rect 1710 48862 1762 48914
rect 16382 48862 16434 48914
rect 16494 48862 16546 48914
rect 20414 48862 20466 48914
rect 20526 48862 20578 48914
rect 22542 48862 22594 48914
rect 22878 48862 22930 48914
rect 22990 48862 23042 48914
rect 26014 48862 26066 48914
rect 27806 48862 27858 48914
rect 31726 48862 31778 48914
rect 2046 48750 2098 48802
rect 2494 48750 2546 48802
rect 9662 48750 9714 48802
rect 12462 48750 12514 48802
rect 14478 48750 14530 48802
rect 14926 48750 14978 48802
rect 16158 48750 16210 48802
rect 18398 48750 18450 48802
rect 18958 48750 19010 48802
rect 19630 48750 19682 48802
rect 20190 48750 20242 48802
rect 22430 48750 22482 48802
rect 23214 48750 23266 48802
rect 27134 48750 27186 48802
rect 37102 48750 37154 48802
rect 38894 48750 38946 48802
rect 19838 48582 19890 48634
rect 19942 48582 19994 48634
rect 20046 48582 20098 48634
rect 50558 48582 50610 48634
rect 50662 48582 50714 48634
rect 50766 48582 50818 48634
rect 3502 48414 3554 48466
rect 16606 48414 16658 48466
rect 22878 48414 22930 48466
rect 30494 48414 30546 48466
rect 31390 48414 31442 48466
rect 39230 48414 39282 48466
rect 7086 48302 7138 48354
rect 7198 48302 7250 48354
rect 10782 48302 10834 48354
rect 19294 48302 19346 48354
rect 19630 48302 19682 48354
rect 21870 48302 21922 48354
rect 23438 48302 23490 48354
rect 23886 48302 23938 48354
rect 23998 48302 24050 48354
rect 26462 48302 26514 48354
rect 27358 48302 27410 48354
rect 29486 48302 29538 48354
rect 30830 48302 30882 48354
rect 31502 48302 31554 48354
rect 31726 48302 31778 48354
rect 38558 48302 38610 48354
rect 39566 48302 39618 48354
rect 6638 48190 6690 48242
rect 9662 48190 9714 48242
rect 10558 48190 10610 48242
rect 11342 48190 11394 48242
rect 11790 48190 11842 48242
rect 14142 48190 14194 48242
rect 15374 48190 15426 48242
rect 18174 48190 18226 48242
rect 18622 48190 18674 48242
rect 20078 48190 20130 48242
rect 21646 48190 21698 48242
rect 22766 48190 22818 48242
rect 23102 48190 23154 48242
rect 23326 48190 23378 48242
rect 23662 48190 23714 48242
rect 24558 48190 24610 48242
rect 26574 48190 26626 48242
rect 27134 48190 27186 48242
rect 29038 48190 29090 48242
rect 29822 48190 29874 48242
rect 31166 48190 31218 48242
rect 33630 48190 33682 48242
rect 4062 48078 4114 48130
rect 6078 48078 6130 48130
rect 10222 48078 10274 48130
rect 14366 48078 14418 48130
rect 15262 48078 15314 48130
rect 16158 48078 16210 48130
rect 17614 48078 17666 48130
rect 18734 48078 18786 48130
rect 20302 48078 20354 48130
rect 22430 48078 22482 48130
rect 32174 48078 32226 48130
rect 33294 48078 33346 48130
rect 7086 47966 7138 48018
rect 11678 47966 11730 48018
rect 13470 47966 13522 48018
rect 13918 47966 13970 48018
rect 15598 47966 15650 48018
rect 16158 47966 16210 48018
rect 16382 47966 16434 48018
rect 17502 47966 17554 48018
rect 23998 47966 24050 48018
rect 4478 47798 4530 47850
rect 4582 47798 4634 47850
rect 4686 47798 4738 47850
rect 35198 47798 35250 47850
rect 35302 47798 35354 47850
rect 35406 47798 35458 47850
rect 3278 47630 3330 47682
rect 16158 47630 16210 47682
rect 16830 47630 16882 47682
rect 18510 47630 18562 47682
rect 19294 47630 19346 47682
rect 2606 47518 2658 47570
rect 7758 47518 7810 47570
rect 16830 47518 16882 47570
rect 18174 47518 18226 47570
rect 32062 47518 32114 47570
rect 32846 47518 32898 47570
rect 34302 47518 34354 47570
rect 35758 47518 35810 47570
rect 37774 47518 37826 47570
rect 39902 47518 39954 47570
rect 2158 47406 2210 47458
rect 3950 47406 4002 47458
rect 6638 47406 6690 47458
rect 7310 47406 7362 47458
rect 8318 47406 8370 47458
rect 8766 47406 8818 47458
rect 10782 47406 10834 47458
rect 12798 47406 12850 47458
rect 13582 47406 13634 47458
rect 13806 47406 13858 47458
rect 14030 47406 14082 47458
rect 14814 47406 14866 47458
rect 15374 47406 15426 47458
rect 15710 47406 15762 47458
rect 16046 47406 16098 47458
rect 17166 47406 17218 47458
rect 18286 47406 18338 47458
rect 19182 47406 19234 47458
rect 19518 47406 19570 47458
rect 19742 47406 19794 47458
rect 20078 47406 20130 47458
rect 25902 47406 25954 47458
rect 27358 47406 27410 47458
rect 29374 47406 29426 47458
rect 30942 47406 30994 47458
rect 31278 47406 31330 47458
rect 33182 47406 33234 47458
rect 33742 47406 33794 47458
rect 34190 47406 34242 47458
rect 34974 47406 35026 47458
rect 35310 47406 35362 47458
rect 38110 47406 38162 47458
rect 39006 47406 39058 47458
rect 42702 47406 42754 47458
rect 3054 47294 3106 47346
rect 4510 47294 4562 47346
rect 6190 47294 6242 47346
rect 9214 47294 9266 47346
rect 12238 47294 12290 47346
rect 17278 47294 17330 47346
rect 18958 47294 19010 47346
rect 26014 47294 26066 47346
rect 28142 47294 28194 47346
rect 29150 47294 29202 47346
rect 33518 47294 33570 47346
rect 34750 47294 34802 47346
rect 42030 47294 42082 47346
rect 3614 47182 3666 47234
rect 12686 47182 12738 47234
rect 14478 47182 14530 47234
rect 16382 47182 16434 47234
rect 17502 47182 17554 47234
rect 18174 47182 18226 47234
rect 20302 47182 20354 47234
rect 20414 47182 20466 47234
rect 24670 47182 24722 47234
rect 26910 47182 26962 47234
rect 34414 47182 34466 47234
rect 35198 47182 35250 47234
rect 38446 47182 38498 47234
rect 39118 47182 39170 47234
rect 39230 47182 39282 47234
rect 39454 47182 39506 47234
rect 19838 47014 19890 47066
rect 19942 47014 19994 47066
rect 20046 47014 20098 47066
rect 50558 47014 50610 47066
rect 50662 47014 50714 47066
rect 50766 47014 50818 47066
rect 2494 46846 2546 46898
rect 13358 46846 13410 46898
rect 16158 46846 16210 46898
rect 33406 46846 33458 46898
rect 38894 46846 38946 46898
rect 40014 46846 40066 46898
rect 40350 46846 40402 46898
rect 41246 46846 41298 46898
rect 1710 46734 1762 46786
rect 2046 46734 2098 46786
rect 2942 46734 2994 46786
rect 3726 46734 3778 46786
rect 4846 46734 4898 46786
rect 6414 46734 6466 46786
rect 7870 46734 7922 46786
rect 10334 46734 10386 46786
rect 11342 46734 11394 46786
rect 13134 46734 13186 46786
rect 19966 46734 20018 46786
rect 27918 46734 27970 46786
rect 33630 46734 33682 46786
rect 36654 46734 36706 46786
rect 39454 46734 39506 46786
rect 40910 46734 40962 46786
rect 41134 46734 41186 46786
rect 41470 46734 41522 46786
rect 3950 46622 4002 46674
rect 4510 46622 4562 46674
rect 6974 46622 7026 46674
rect 7310 46622 7362 46674
rect 10446 46622 10498 46674
rect 11454 46622 11506 46674
rect 13582 46622 13634 46674
rect 14142 46622 14194 46674
rect 14702 46622 14754 46674
rect 15038 46622 15090 46674
rect 20302 46622 20354 46674
rect 25230 46622 25282 46674
rect 32622 46622 32674 46674
rect 33070 46622 33122 46674
rect 33294 46622 33346 46674
rect 37326 46622 37378 46674
rect 39118 46622 39170 46674
rect 3838 46510 3890 46562
rect 5966 46510 6018 46562
rect 15710 46510 15762 46562
rect 22766 46510 22818 46562
rect 24334 46510 24386 46562
rect 24782 46510 24834 46562
rect 34526 46510 34578 46562
rect 3054 46398 3106 46450
rect 15038 46398 15090 46450
rect 20302 46398 20354 46450
rect 4478 46230 4530 46282
rect 4582 46230 4634 46282
rect 4686 46230 4738 46282
rect 35198 46230 35250 46282
rect 35302 46230 35354 46282
rect 35406 46230 35458 46282
rect 14702 46062 14754 46114
rect 15038 46062 15090 46114
rect 7310 45950 7362 46002
rect 9886 45950 9938 46002
rect 14478 45950 14530 46002
rect 15038 45950 15090 46002
rect 22206 45950 22258 46002
rect 22654 45950 22706 46002
rect 27806 45950 27858 46002
rect 32062 45950 32114 46002
rect 32846 45950 32898 46002
rect 33742 45950 33794 46002
rect 34750 45950 34802 46002
rect 41022 45950 41074 46002
rect 3950 45838 4002 45890
rect 6862 45838 6914 45890
rect 7646 45838 7698 45890
rect 8654 45838 8706 45890
rect 10334 45838 10386 45890
rect 12126 45838 12178 45890
rect 13918 45838 13970 45890
rect 16046 45838 16098 45890
rect 16494 45838 16546 45890
rect 16718 45838 16770 45890
rect 19966 45838 20018 45890
rect 20078 45838 20130 45890
rect 21646 45838 21698 45890
rect 21982 45838 22034 45890
rect 24446 45838 24498 45890
rect 24782 45838 24834 45890
rect 26798 45838 26850 45890
rect 29374 45838 29426 45890
rect 31838 45838 31890 45890
rect 32734 45838 32786 45890
rect 32958 45838 33010 45890
rect 33406 45838 33458 45890
rect 34190 45838 34242 45890
rect 34638 45838 34690 45890
rect 34862 45838 34914 45890
rect 38558 45838 38610 45890
rect 38670 45838 38722 45890
rect 41582 45838 41634 45890
rect 41918 45838 41970 45890
rect 1710 45726 1762 45778
rect 4510 45726 4562 45778
rect 6526 45726 6578 45778
rect 9326 45726 9378 45778
rect 10894 45726 10946 45778
rect 16270 45726 16322 45778
rect 17838 45726 17890 45778
rect 23662 45726 23714 45778
rect 24222 45726 24274 45778
rect 24558 45726 24610 45778
rect 24894 45726 24946 45778
rect 27358 45726 27410 45778
rect 29486 45726 29538 45778
rect 31726 45726 31778 45778
rect 41358 45726 41410 45778
rect 2046 45614 2098 45666
rect 2494 45614 2546 45666
rect 6638 45614 6690 45666
rect 8094 45614 8146 45666
rect 10446 45614 10498 45666
rect 16158 45614 16210 45666
rect 17390 45614 17442 45666
rect 19742 45614 19794 45666
rect 20638 45614 20690 45666
rect 21422 45614 21474 45666
rect 21534 45614 21586 45666
rect 22430 45614 22482 45666
rect 23102 45614 23154 45666
rect 41806 45614 41858 45666
rect 19838 45446 19890 45498
rect 19942 45446 19994 45498
rect 20046 45446 20098 45498
rect 50558 45446 50610 45498
rect 50662 45446 50714 45498
rect 50766 45446 50818 45498
rect 2606 45278 2658 45330
rect 3166 45278 3218 45330
rect 8206 45278 8258 45330
rect 19070 45278 19122 45330
rect 21422 45278 21474 45330
rect 22654 45278 22706 45330
rect 23438 45278 23490 45330
rect 25678 45278 25730 45330
rect 27582 45278 27634 45330
rect 32510 45278 32562 45330
rect 40238 45278 40290 45330
rect 7982 45166 8034 45218
rect 10222 45166 10274 45218
rect 19406 45166 19458 45218
rect 19630 45166 19682 45218
rect 21646 45166 21698 45218
rect 22542 45166 22594 45218
rect 25902 45166 25954 45218
rect 26238 45166 26290 45218
rect 28702 45166 28754 45218
rect 33182 45166 33234 45218
rect 33406 45166 33458 45218
rect 42366 45166 42418 45218
rect 2494 45054 2546 45106
rect 2830 45054 2882 45106
rect 3054 45054 3106 45106
rect 4174 45054 4226 45106
rect 6862 45054 6914 45106
rect 6974 45054 7026 45106
rect 7758 45054 7810 45106
rect 11118 45054 11170 45106
rect 11454 45054 11506 45106
rect 13806 45054 13858 45106
rect 19966 45054 20018 45106
rect 20750 45054 20802 45106
rect 21870 45054 21922 45106
rect 22318 45054 22370 45106
rect 22878 45054 22930 45106
rect 25566 45054 25618 45106
rect 26126 45054 26178 45106
rect 29934 45054 29986 45106
rect 33854 45054 33906 45106
rect 39678 45054 39730 45106
rect 40126 45054 40178 45106
rect 40350 45054 40402 45106
rect 41582 45054 41634 45106
rect 3838 44942 3890 44994
rect 6750 44942 6802 44994
rect 8206 44942 8258 44994
rect 11566 44942 11618 44994
rect 14366 44942 14418 44994
rect 18622 44942 18674 44994
rect 20302 44942 20354 44994
rect 24334 44942 24386 44994
rect 24670 44942 24722 44994
rect 36990 44942 37042 44994
rect 44494 44942 44546 44994
rect 3166 44830 3218 44882
rect 20526 44830 20578 44882
rect 20974 44830 21026 44882
rect 22094 44830 22146 44882
rect 23102 44830 23154 44882
rect 33518 44830 33570 44882
rect 4478 44662 4530 44714
rect 4582 44662 4634 44714
rect 4686 44662 4738 44714
rect 35198 44662 35250 44714
rect 35302 44662 35354 44714
rect 35406 44662 35458 44714
rect 22094 44494 22146 44546
rect 25790 44494 25842 44546
rect 27134 44494 27186 44546
rect 34414 44494 34466 44546
rect 8542 44382 8594 44434
rect 13806 44382 13858 44434
rect 14814 44382 14866 44434
rect 16158 44382 16210 44434
rect 23438 44382 23490 44434
rect 24670 44382 24722 44434
rect 26126 44382 26178 44434
rect 28478 44382 28530 44434
rect 29374 44382 29426 44434
rect 35422 44382 35474 44434
rect 37550 44382 37602 44434
rect 38558 44382 38610 44434
rect 6862 44270 6914 44322
rect 10222 44270 10274 44322
rect 10446 44270 10498 44322
rect 11006 44270 11058 44322
rect 11230 44270 11282 44322
rect 11454 44270 11506 44322
rect 14254 44270 14306 44322
rect 15262 44270 15314 44322
rect 15710 44270 15762 44322
rect 16382 44270 16434 44322
rect 16606 44270 16658 44322
rect 16830 44270 16882 44322
rect 17502 44270 17554 44322
rect 20750 44270 20802 44322
rect 21310 44270 21362 44322
rect 21646 44270 21698 44322
rect 22990 44270 23042 44322
rect 24446 44270 24498 44322
rect 26350 44270 26402 44322
rect 26686 44270 26738 44322
rect 29598 44270 29650 44322
rect 30830 44270 30882 44322
rect 33294 44270 33346 44322
rect 34190 44270 34242 44322
rect 34750 44270 34802 44322
rect 39006 44270 39058 44322
rect 39118 44270 39170 44322
rect 39566 44270 39618 44322
rect 5742 44158 5794 44210
rect 8094 44158 8146 44210
rect 10558 44158 10610 44210
rect 17390 44158 17442 44210
rect 19182 44158 19234 44210
rect 19854 44158 19906 44210
rect 21534 44158 21586 44210
rect 22654 44158 22706 44210
rect 24222 44158 24274 44210
rect 26462 44158 26514 44210
rect 29934 44158 29986 44210
rect 30606 44158 30658 44210
rect 32958 44158 33010 44210
rect 34974 44158 35026 44210
rect 37438 44158 37490 44210
rect 12238 44046 12290 44098
rect 17278 44046 17330 44098
rect 25006 44046 25058 44098
rect 27470 44046 27522 44098
rect 27806 44046 27858 44098
rect 32622 44046 32674 44098
rect 34638 44046 34690 44098
rect 39342 44046 39394 44098
rect 19838 43878 19890 43930
rect 19942 43878 19994 43930
rect 20046 43878 20098 43930
rect 50558 43878 50610 43930
rect 50662 43878 50714 43930
rect 50766 43878 50818 43930
rect 7198 43710 7250 43762
rect 13246 43710 13298 43762
rect 17502 43710 17554 43762
rect 22318 43710 22370 43762
rect 23774 43710 23826 43762
rect 28254 43710 28306 43762
rect 2270 43598 2322 43650
rect 2718 43598 2770 43650
rect 5294 43598 5346 43650
rect 6526 43598 6578 43650
rect 7758 43598 7810 43650
rect 11006 43598 11058 43650
rect 13134 43598 13186 43650
rect 17390 43598 17442 43650
rect 17614 43598 17666 43650
rect 18734 43598 18786 43650
rect 21758 43598 21810 43650
rect 24558 43598 24610 43650
rect 25342 43598 25394 43650
rect 26238 43598 26290 43650
rect 26574 43598 26626 43650
rect 29150 43598 29202 43650
rect 31502 43598 31554 43650
rect 31726 43598 31778 43650
rect 32062 43598 32114 43650
rect 32622 43598 32674 43650
rect 33070 43598 33122 43650
rect 33406 43598 33458 43650
rect 34638 43598 34690 43650
rect 39342 43598 39394 43650
rect 41246 43598 41298 43650
rect 2494 43486 2546 43538
rect 2942 43486 2994 43538
rect 3502 43486 3554 43538
rect 4846 43486 4898 43538
rect 6862 43486 6914 43538
rect 10110 43486 10162 43538
rect 12798 43486 12850 43538
rect 13470 43486 13522 43538
rect 13918 43486 13970 43538
rect 17838 43486 17890 43538
rect 18174 43486 18226 43538
rect 18622 43486 18674 43538
rect 20638 43486 20690 43538
rect 23438 43486 23490 43538
rect 24222 43486 24274 43538
rect 25566 43486 25618 43538
rect 25790 43486 25842 43538
rect 28142 43486 28194 43538
rect 28590 43486 28642 43538
rect 33966 43486 34018 43538
rect 40014 43486 40066 43538
rect 41134 43486 41186 43538
rect 41358 43486 41410 43538
rect 41694 43486 41746 43538
rect 1822 43374 1874 43426
rect 2830 43374 2882 43426
rect 4062 43374 4114 43426
rect 4510 43374 4562 43426
rect 5854 43374 5906 43426
rect 9998 43374 10050 43426
rect 11342 43374 11394 43426
rect 12462 43374 12514 43426
rect 14478 43374 14530 43426
rect 23102 43374 23154 43426
rect 25230 43374 25282 43426
rect 36766 43374 36818 43426
rect 37214 43374 37266 43426
rect 6862 43262 6914 43314
rect 9662 43262 9714 43314
rect 9774 43262 9826 43314
rect 11454 43262 11506 43314
rect 24670 43262 24722 43314
rect 4478 43094 4530 43146
rect 4582 43094 4634 43146
rect 4686 43094 4738 43146
rect 35198 43094 35250 43146
rect 35302 43094 35354 43146
rect 35406 43094 35458 43146
rect 8318 42926 8370 42978
rect 22654 42926 22706 42978
rect 23438 42926 23490 42978
rect 23998 42926 24050 42978
rect 25006 42926 25058 42978
rect 30046 42926 30098 42978
rect 7982 42814 8034 42866
rect 13918 42814 13970 42866
rect 21758 42814 21810 42866
rect 23662 42814 23714 42866
rect 38670 42814 38722 42866
rect 39118 42814 39170 42866
rect 44046 42814 44098 42866
rect 1822 42702 1874 42754
rect 7870 42702 7922 42754
rect 8206 42702 8258 42754
rect 8766 42702 8818 42754
rect 10782 42702 10834 42754
rect 13470 42702 13522 42754
rect 17614 42702 17666 42754
rect 18062 42702 18114 42754
rect 24446 42702 24498 42754
rect 24670 42702 24722 42754
rect 25566 42702 25618 42754
rect 27806 42702 27858 42754
rect 29374 42702 29426 42754
rect 29934 42702 29986 42754
rect 30270 42702 30322 42754
rect 31054 42702 31106 42754
rect 33518 42702 33570 42754
rect 38558 42702 38610 42754
rect 39230 42702 39282 42754
rect 40126 42702 40178 42754
rect 40798 42702 40850 42754
rect 41134 42702 41186 42754
rect 2046 42590 2098 42642
rect 2718 42590 2770 42642
rect 2830 42590 2882 42642
rect 8878 42590 8930 42642
rect 11902 42590 11954 42642
rect 23886 42590 23938 42642
rect 25454 42590 25506 42642
rect 27358 42590 27410 42642
rect 30830 42590 30882 42642
rect 32958 42590 33010 42642
rect 39006 42590 39058 42642
rect 39454 42590 39506 42642
rect 40574 42590 40626 42642
rect 41918 42590 41970 42642
rect 3054 42478 3106 42530
rect 10334 42478 10386 42530
rect 20750 42478 20802 42530
rect 21310 42478 21362 42530
rect 22654 42478 22706 42530
rect 23214 42478 23266 42530
rect 23998 42478 24050 42530
rect 28366 42478 28418 42530
rect 32846 42478 32898 42530
rect 34638 42478 34690 42530
rect 40462 42478 40514 42530
rect 19838 42310 19890 42362
rect 19942 42310 19994 42362
rect 20046 42310 20098 42362
rect 50558 42310 50610 42362
rect 50662 42310 50714 42362
rect 50766 42310 50818 42362
rect 3502 42142 3554 42194
rect 8878 42142 8930 42194
rect 16718 42142 16770 42194
rect 23662 42142 23714 42194
rect 29374 42142 29426 42194
rect 35422 42142 35474 42194
rect 2270 42030 2322 42082
rect 6414 42030 6466 42082
rect 8990 42030 9042 42082
rect 11118 42030 11170 42082
rect 12126 42030 12178 42082
rect 17838 42030 17890 42082
rect 17950 42030 18002 42082
rect 27918 42030 27970 42082
rect 30494 42030 30546 42082
rect 34526 42030 34578 42082
rect 34974 42030 35026 42082
rect 35198 42030 35250 42082
rect 41022 42030 41074 42082
rect 2494 41918 2546 41970
rect 2718 41918 2770 41970
rect 2830 41918 2882 41970
rect 5294 41918 5346 41970
rect 7422 41918 7474 41970
rect 11454 41918 11506 41970
rect 12238 41918 12290 41970
rect 16606 41918 16658 41970
rect 18174 41918 18226 41970
rect 18622 41918 18674 41970
rect 20190 41918 20242 41970
rect 20414 41918 20466 41970
rect 20638 41918 20690 41970
rect 20862 41918 20914 41970
rect 20974 41918 21026 41970
rect 22094 41918 22146 41970
rect 22206 41918 22258 41970
rect 22430 41918 22482 41970
rect 22878 41918 22930 41970
rect 29598 41918 29650 41970
rect 29934 41918 29986 41970
rect 33518 41918 33570 41970
rect 35758 41918 35810 41970
rect 1822 41806 1874 41858
rect 2606 41806 2658 41858
rect 4062 41806 4114 41858
rect 13022 41806 13074 41858
rect 19854 41806 19906 41858
rect 21534 41806 21586 41858
rect 21870 41806 21922 41858
rect 23214 41806 23266 41858
rect 24670 41806 24722 41858
rect 25342 41806 25394 41858
rect 26574 41806 26626 41858
rect 27246 41806 27298 41858
rect 34078 41806 34130 41858
rect 36206 41806 36258 41858
rect 39902 41806 39954 41858
rect 16718 41694 16770 41746
rect 18510 41694 18562 41746
rect 18846 41694 18898 41746
rect 18958 41694 19010 41746
rect 34302 41694 34354 41746
rect 34638 41694 34690 41746
rect 35422 41694 35474 41746
rect 40910 41694 40962 41746
rect 4478 41526 4530 41578
rect 4582 41526 4634 41578
rect 4686 41526 4738 41578
rect 35198 41526 35250 41578
rect 35302 41526 35354 41578
rect 35406 41526 35458 41578
rect 13806 41358 13858 41410
rect 14254 41358 14306 41410
rect 21758 41358 21810 41410
rect 22094 41358 22146 41410
rect 28254 41358 28306 41410
rect 30046 41358 30098 41410
rect 35310 41358 35362 41410
rect 7646 41246 7698 41298
rect 9550 41246 9602 41298
rect 12574 41246 12626 41298
rect 18398 41246 18450 41298
rect 24558 41246 24610 41298
rect 27918 41246 27970 41298
rect 35982 41246 36034 41298
rect 1710 41134 1762 41186
rect 5854 41134 5906 41186
rect 9102 41134 9154 41186
rect 9326 41134 9378 41186
rect 10334 41134 10386 41186
rect 10894 41134 10946 41186
rect 11902 41134 11954 41186
rect 14030 41134 14082 41186
rect 17166 41134 17218 41186
rect 17614 41134 17666 41186
rect 19630 41134 19682 41186
rect 19966 41134 20018 41186
rect 20862 41134 20914 41186
rect 21422 41134 21474 41186
rect 21534 41134 21586 41186
rect 21982 41134 22034 41186
rect 23326 41134 23378 41186
rect 24894 41134 24946 41186
rect 26910 41134 26962 41186
rect 27134 41134 27186 41186
rect 28366 41134 28418 41186
rect 29150 41134 29202 41186
rect 29374 41134 29426 41186
rect 29598 41134 29650 41186
rect 31278 41134 31330 41186
rect 32958 41134 33010 41186
rect 33518 41134 33570 41186
rect 34750 41134 34802 41186
rect 35310 41134 35362 41186
rect 2046 41022 2098 41074
rect 2382 41022 2434 41074
rect 2718 41022 2770 41074
rect 6414 41022 6466 41074
rect 12126 41022 12178 41074
rect 13582 41022 13634 41074
rect 15710 41022 15762 41074
rect 18734 41022 18786 41074
rect 19854 41022 19906 41074
rect 20526 41022 20578 41074
rect 23886 41022 23938 41074
rect 25118 41022 25170 41074
rect 31054 41022 31106 41074
rect 34974 41022 35026 41074
rect 35870 41022 35922 41074
rect 7870 40910 7922 40962
rect 9550 40910 9602 40962
rect 14702 40910 14754 40962
rect 15038 40910 15090 40962
rect 20638 40910 20690 40962
rect 22542 40910 22594 40962
rect 22990 40910 23042 40962
rect 30382 40910 30434 40962
rect 33070 40910 33122 40962
rect 35198 40910 35250 40962
rect 36094 40910 36146 40962
rect 19838 40742 19890 40794
rect 19942 40742 19994 40794
rect 20046 40742 20098 40794
rect 50558 40742 50610 40794
rect 50662 40742 50714 40794
rect 50766 40742 50818 40794
rect 12238 40574 12290 40626
rect 13022 40574 13074 40626
rect 16382 40574 16434 40626
rect 18174 40574 18226 40626
rect 19518 40574 19570 40626
rect 21086 40574 21138 40626
rect 24110 40574 24162 40626
rect 26686 40574 26738 40626
rect 27358 40574 27410 40626
rect 27694 40574 27746 40626
rect 34078 40574 34130 40626
rect 34526 40574 34578 40626
rect 35758 40574 35810 40626
rect 36318 40574 36370 40626
rect 2046 40462 2098 40514
rect 4174 40462 4226 40514
rect 6190 40462 6242 40514
rect 9662 40462 9714 40514
rect 11678 40462 11730 40514
rect 15934 40462 15986 40514
rect 16158 40462 16210 40514
rect 17726 40462 17778 40514
rect 18734 40462 18786 40514
rect 25230 40462 25282 40514
rect 34974 40462 35026 40514
rect 37774 40462 37826 40514
rect 1710 40350 1762 40402
rect 2494 40350 2546 40402
rect 3390 40350 3442 40402
rect 3614 40350 3666 40402
rect 5742 40350 5794 40402
rect 8094 40350 8146 40402
rect 8430 40350 8482 40402
rect 9102 40350 9154 40402
rect 9886 40350 9938 40402
rect 11454 40350 11506 40402
rect 12798 40350 12850 40402
rect 13358 40350 13410 40402
rect 14366 40350 14418 40402
rect 15374 40350 15426 40402
rect 16606 40350 16658 40402
rect 17502 40350 17554 40402
rect 18846 40350 18898 40402
rect 19070 40350 19122 40402
rect 22542 40350 22594 40402
rect 28590 40350 28642 40402
rect 28814 40350 28866 40402
rect 30158 40350 30210 40402
rect 30830 40350 30882 40402
rect 31390 40350 31442 40402
rect 35310 40350 35362 40402
rect 35422 40350 35474 40402
rect 35534 40350 35586 40402
rect 36990 40350 37042 40402
rect 5406 40238 5458 40290
rect 8766 40238 8818 40290
rect 11902 40238 11954 40290
rect 12910 40238 12962 40290
rect 14814 40238 14866 40290
rect 18510 40238 18562 40290
rect 26126 40238 26178 40290
rect 30382 40238 30434 40290
rect 34638 40238 34690 40290
rect 39902 40238 39954 40290
rect 25342 40126 25394 40178
rect 25566 40126 25618 40178
rect 25678 40126 25730 40178
rect 26350 40126 26402 40178
rect 34302 40126 34354 40178
rect 4478 39958 4530 40010
rect 4582 39958 4634 40010
rect 4686 39958 4738 40010
rect 35198 39958 35250 40010
rect 35302 39958 35354 40010
rect 35406 39958 35458 40010
rect 27918 39790 27970 39842
rect 28030 39790 28082 39842
rect 28254 39790 28306 39842
rect 30270 39790 30322 39842
rect 8094 39678 8146 39730
rect 11118 39678 11170 39730
rect 20078 39678 20130 39730
rect 22094 39678 22146 39730
rect 26462 39678 26514 39730
rect 27582 39678 27634 39730
rect 29486 39678 29538 39730
rect 32174 39678 32226 39730
rect 3950 39566 4002 39618
rect 5070 39566 5122 39618
rect 6750 39566 6802 39618
rect 7982 39566 8034 39618
rect 10558 39566 10610 39618
rect 10782 39566 10834 39618
rect 15038 39566 15090 39618
rect 16382 39566 16434 39618
rect 17390 39566 17442 39618
rect 18958 39566 19010 39618
rect 21310 39566 21362 39618
rect 23326 39566 23378 39618
rect 27022 39566 27074 39618
rect 28478 39566 28530 39618
rect 30046 39566 30098 39618
rect 30606 39566 30658 39618
rect 30830 39566 30882 39618
rect 31502 39566 31554 39618
rect 31726 39566 31778 39618
rect 33966 39566 34018 39618
rect 34302 39566 34354 39618
rect 2830 39454 2882 39506
rect 3054 39454 3106 39506
rect 3390 39454 3442 39506
rect 4958 39454 5010 39506
rect 7198 39454 7250 39506
rect 8206 39454 8258 39506
rect 14702 39454 14754 39506
rect 18174 39454 18226 39506
rect 23886 39454 23938 39506
rect 27134 39454 27186 39506
rect 33742 39454 33794 39506
rect 34638 39454 34690 39506
rect 2942 39342 2994 39394
rect 3502 39342 3554 39394
rect 6078 39342 6130 39394
rect 11006 39342 11058 39394
rect 14142 39342 14194 39394
rect 15150 39342 15202 39394
rect 19518 39342 19570 39394
rect 22990 39342 23042 39394
rect 19838 39174 19890 39226
rect 19942 39174 19994 39226
rect 20046 39174 20098 39226
rect 50558 39174 50610 39226
rect 50662 39174 50714 39226
rect 50766 39174 50818 39226
rect 5294 39006 5346 39058
rect 5854 39006 5906 39058
rect 11790 39006 11842 39058
rect 13022 39006 13074 39058
rect 15038 39006 15090 39058
rect 15262 39006 15314 39058
rect 19406 39006 19458 39058
rect 22206 39006 22258 39058
rect 25118 39006 25170 39058
rect 27582 39006 27634 39058
rect 28702 39006 28754 39058
rect 29262 39006 29314 39058
rect 2382 38894 2434 38946
rect 3502 38894 3554 38946
rect 5742 38894 5794 38946
rect 7310 38894 7362 38946
rect 21310 38894 21362 38946
rect 24222 38894 24274 38946
rect 26686 38894 26738 38946
rect 27918 38894 27970 38946
rect 30942 38894 30994 38946
rect 32398 38894 32450 38946
rect 34414 38894 34466 38946
rect 35310 38894 35362 38946
rect 38222 38894 38274 38946
rect 2606 38782 2658 38834
rect 3838 38782 3890 38834
rect 4286 38782 4338 38834
rect 5630 38782 5682 38834
rect 6750 38782 6802 38834
rect 7758 38782 7810 38834
rect 7982 38782 8034 38834
rect 12350 38782 12402 38834
rect 12798 38782 12850 38834
rect 13918 38782 13970 38834
rect 14478 38782 14530 38834
rect 14814 38782 14866 38834
rect 15486 38782 15538 38834
rect 21198 38782 21250 38834
rect 21534 38782 21586 38834
rect 21982 38782 22034 38834
rect 23774 38782 23826 38834
rect 24670 38782 24722 38834
rect 25790 38782 25842 38834
rect 26014 38782 26066 38834
rect 26910 38782 26962 38834
rect 27134 38782 27186 38834
rect 31166 38782 31218 38834
rect 31726 38782 31778 38834
rect 32510 38782 32562 38834
rect 34302 38782 34354 38834
rect 36766 38782 36818 38834
rect 37438 38782 37490 38834
rect 1822 38670 1874 38722
rect 8094 38670 8146 38722
rect 8654 38670 8706 38722
rect 16270 38670 16322 38722
rect 18062 38670 18114 38722
rect 18622 38670 18674 38722
rect 19070 38670 19122 38722
rect 20302 38670 20354 38722
rect 20974 38670 21026 38722
rect 22766 38670 22818 38722
rect 23214 38670 23266 38722
rect 7646 38558 7698 38610
rect 15374 38558 15426 38610
rect 23998 38558 24050 38610
rect 24558 38670 24610 38722
rect 25566 38670 25618 38722
rect 26238 38670 26290 38722
rect 26574 38670 26626 38722
rect 33630 38670 33682 38722
rect 40350 38670 40402 38722
rect 4478 38390 4530 38442
rect 4582 38390 4634 38442
rect 4686 38390 4738 38442
rect 35198 38390 35250 38442
rect 35302 38390 35354 38442
rect 35406 38390 35458 38442
rect 4958 38222 5010 38274
rect 11230 38222 11282 38274
rect 3950 38110 4002 38162
rect 7422 38110 7474 38162
rect 12238 38110 12290 38162
rect 13358 38110 13410 38162
rect 15150 38110 15202 38162
rect 2494 37998 2546 38050
rect 3054 37998 3106 38050
rect 3614 37998 3666 38050
rect 4734 37998 4786 38050
rect 5630 37998 5682 38050
rect 6526 37998 6578 38050
rect 7534 37998 7586 38050
rect 9214 37998 9266 38050
rect 9550 37998 9602 38050
rect 9998 37998 10050 38050
rect 11790 37998 11842 38050
rect 11902 37998 11954 38050
rect 12350 37998 12402 38050
rect 14030 37998 14082 38050
rect 15038 37998 15090 38050
rect 15598 37998 15650 38050
rect 1710 37886 1762 37938
rect 2606 37886 2658 37938
rect 4062 37886 4114 37938
rect 4286 37886 4338 37938
rect 6750 37886 6802 37938
rect 10894 37886 10946 37938
rect 11342 37886 11394 37938
rect 13470 37886 13522 37938
rect 14478 37886 14530 37938
rect 15934 37886 15986 37938
rect 16606 38222 16658 38274
rect 19070 38222 19122 38274
rect 20638 38222 20690 38274
rect 37774 38222 37826 38274
rect 19630 38110 19682 38162
rect 22878 38110 22930 38162
rect 26238 38110 26290 38162
rect 28366 38110 28418 38162
rect 30046 38110 30098 38162
rect 32846 38110 32898 38162
rect 34190 38110 34242 38162
rect 36430 38110 36482 38162
rect 37214 38110 37266 38162
rect 17166 37998 17218 38050
rect 17838 37998 17890 38050
rect 18286 37998 18338 38050
rect 18510 37998 18562 38050
rect 18734 37998 18786 38050
rect 18958 37998 19010 38050
rect 19966 37998 20018 38050
rect 20302 37998 20354 38050
rect 24110 37998 24162 38050
rect 26126 37998 26178 38050
rect 28590 37998 28642 38050
rect 29822 37998 29874 38050
rect 30494 37998 30546 38050
rect 31838 37998 31890 38050
rect 33294 37998 33346 38050
rect 37998 37998 38050 38050
rect 38222 37998 38274 38050
rect 38446 37998 38498 38050
rect 17726 37886 17778 37938
rect 19742 37886 19794 37938
rect 24222 37886 24274 37938
rect 27246 37886 27298 37938
rect 28254 37886 28306 37938
rect 30606 37886 30658 37938
rect 32062 37886 32114 37938
rect 32174 37886 32226 37938
rect 2046 37774 2098 37826
rect 2830 37774 2882 37826
rect 6190 37774 6242 37826
rect 6862 37774 6914 37826
rect 10670 37774 10722 37826
rect 11118 37774 11170 37826
rect 12126 37774 12178 37826
rect 12798 37774 12850 37826
rect 13694 37774 13746 37826
rect 13918 37774 13970 37826
rect 15710 37774 15762 37826
rect 16382 37774 16434 37826
rect 17278 37774 17330 37826
rect 17502 37774 17554 37826
rect 21534 37774 21586 37826
rect 21982 37774 22034 37826
rect 22542 37774 22594 37826
rect 23438 37774 23490 37826
rect 23774 37774 23826 37826
rect 29710 37774 29762 37826
rect 33742 37774 33794 37826
rect 19838 37606 19890 37658
rect 19942 37606 19994 37658
rect 20046 37606 20098 37658
rect 50558 37606 50610 37658
rect 50662 37606 50714 37658
rect 50766 37606 50818 37658
rect 2606 37438 2658 37490
rect 2830 37438 2882 37490
rect 6302 37438 6354 37490
rect 8206 37438 8258 37490
rect 10558 37438 10610 37490
rect 12574 37438 12626 37490
rect 13022 37438 13074 37490
rect 18622 37438 18674 37490
rect 19182 37438 19234 37490
rect 19406 37438 19458 37490
rect 25230 37438 25282 37490
rect 26014 37438 26066 37490
rect 26798 37438 26850 37490
rect 29598 37438 29650 37490
rect 29710 37438 29762 37490
rect 32062 37438 32114 37490
rect 39902 37438 39954 37490
rect 2046 37326 2098 37378
rect 2494 37326 2546 37378
rect 9774 37326 9826 37378
rect 12126 37326 12178 37378
rect 15822 37326 15874 37378
rect 16494 37326 16546 37378
rect 17838 37326 17890 37378
rect 18286 37326 18338 37378
rect 18398 37326 18450 37378
rect 21198 37326 21250 37378
rect 25454 37326 25506 37378
rect 25566 37326 25618 37378
rect 26238 37326 26290 37378
rect 29038 37326 29090 37378
rect 29486 37326 29538 37378
rect 35870 37326 35922 37378
rect 39566 37326 39618 37378
rect 40238 37326 40290 37378
rect 1710 37214 1762 37266
rect 7758 37214 7810 37266
rect 8654 37214 8706 37266
rect 8766 37214 8818 37266
rect 8990 37214 9042 37266
rect 9662 37214 9714 37266
rect 9886 37214 9938 37266
rect 10110 37214 10162 37266
rect 11902 37214 11954 37266
rect 15150 37214 15202 37266
rect 15374 37214 15426 37266
rect 16046 37214 16098 37266
rect 16270 37214 16322 37266
rect 17502 37214 17554 37266
rect 19070 37214 19122 37266
rect 20078 37214 20130 37266
rect 22654 37214 22706 37266
rect 22878 37214 22930 37266
rect 23214 37214 23266 37266
rect 23550 37214 23602 37266
rect 26574 37214 26626 37266
rect 27694 37214 27746 37266
rect 29822 37214 29874 37266
rect 30046 37214 30098 37266
rect 31054 37214 31106 37266
rect 31278 37214 31330 37266
rect 31502 37214 31554 37266
rect 32286 37214 32338 37266
rect 34190 37214 34242 37266
rect 34750 37214 34802 37266
rect 35086 37214 35138 37266
rect 38670 37214 38722 37266
rect 3166 37102 3218 37154
rect 7422 37102 7474 37154
rect 14926 37102 14978 37154
rect 16158 37102 16210 37154
rect 21422 37102 21474 37154
rect 27246 37102 27298 37154
rect 27918 37102 27970 37154
rect 28478 37102 28530 37154
rect 31950 37102 32002 37154
rect 37998 37102 38050 37154
rect 39118 37102 39170 37154
rect 27470 36990 27522 37042
rect 30494 36990 30546 37042
rect 40350 36990 40402 37042
rect 4478 36822 4530 36874
rect 4582 36822 4634 36874
rect 4686 36822 4738 36874
rect 35198 36822 35250 36874
rect 35302 36822 35354 36874
rect 35406 36822 35458 36874
rect 14142 36654 14194 36706
rect 3614 36542 3666 36594
rect 7086 36542 7138 36594
rect 7982 36542 8034 36594
rect 8206 36542 8258 36594
rect 12910 36542 12962 36594
rect 18062 36542 18114 36594
rect 19294 36542 19346 36594
rect 19854 36542 19906 36594
rect 27582 36542 27634 36594
rect 31726 36542 31778 36594
rect 37326 36542 37378 36594
rect 39342 36542 39394 36594
rect 2494 36430 2546 36482
rect 2718 36430 2770 36482
rect 3278 36430 3330 36482
rect 5742 36430 5794 36482
rect 8654 36430 8706 36482
rect 14366 36430 14418 36482
rect 20414 36430 20466 36482
rect 20750 36430 20802 36482
rect 22542 36430 22594 36482
rect 24222 36430 24274 36482
rect 25342 36430 25394 36482
rect 25790 36430 25842 36482
rect 26014 36430 26066 36482
rect 28702 36430 28754 36482
rect 32734 36430 32786 36482
rect 33182 36430 33234 36482
rect 34414 36430 34466 36482
rect 36206 36430 36258 36482
rect 37998 36430 38050 36482
rect 38558 36430 38610 36482
rect 1934 36318 1986 36370
rect 3838 36318 3890 36370
rect 5966 36318 6018 36370
rect 6750 36318 6802 36370
rect 13806 36318 13858 36370
rect 17502 36318 17554 36370
rect 18062 36318 18114 36370
rect 18286 36318 18338 36370
rect 22990 36318 23042 36370
rect 28366 36318 28418 36370
rect 35646 36318 35698 36370
rect 4286 36206 4338 36258
rect 4846 36206 4898 36258
rect 8990 36206 9042 36258
rect 10558 36206 10610 36258
rect 14030 36206 14082 36258
rect 17838 36206 17890 36258
rect 18958 36206 19010 36258
rect 20302 36206 20354 36258
rect 20638 36206 20690 36258
rect 21534 36206 21586 36258
rect 21870 36206 21922 36258
rect 23886 36206 23938 36258
rect 28030 36206 28082 36258
rect 28478 36206 28530 36258
rect 29262 36206 29314 36258
rect 29710 36206 29762 36258
rect 32286 36206 32338 36258
rect 33854 36206 33906 36258
rect 40126 36206 40178 36258
rect 40910 36206 40962 36258
rect 19838 36038 19890 36090
rect 19942 36038 19994 36090
rect 20046 36038 20098 36090
rect 50558 36038 50610 36090
rect 50662 36038 50714 36090
rect 50766 36038 50818 36090
rect 2494 35870 2546 35922
rect 3502 35870 3554 35922
rect 4622 35870 4674 35922
rect 5742 35870 5794 35922
rect 7646 35870 7698 35922
rect 10110 35870 10162 35922
rect 10446 35870 10498 35922
rect 12014 35870 12066 35922
rect 12574 35870 12626 35922
rect 15038 35870 15090 35922
rect 19070 35870 19122 35922
rect 19742 35870 19794 35922
rect 20862 35870 20914 35922
rect 27470 35870 27522 35922
rect 28254 35870 28306 35922
rect 28478 35870 28530 35922
rect 33406 35870 33458 35922
rect 40350 35870 40402 35922
rect 40910 35870 40962 35922
rect 2270 35758 2322 35810
rect 3726 35758 3778 35810
rect 10334 35758 10386 35810
rect 14814 35758 14866 35810
rect 17726 35758 17778 35810
rect 19294 35758 19346 35810
rect 19966 35758 20018 35810
rect 20526 35758 20578 35810
rect 22878 35758 22930 35810
rect 23886 35758 23938 35810
rect 25454 35758 25506 35810
rect 33854 35758 33906 35810
rect 36430 35758 36482 35810
rect 37438 35758 37490 35810
rect 37662 35758 37714 35810
rect 39230 35758 39282 35810
rect 2606 35646 2658 35698
rect 2718 35646 2770 35698
rect 2830 35646 2882 35698
rect 3166 35646 3218 35698
rect 9774 35646 9826 35698
rect 12126 35646 12178 35698
rect 13918 35646 13970 35698
rect 14702 35646 14754 35698
rect 17614 35646 17666 35698
rect 18734 35646 18786 35698
rect 20078 35646 20130 35698
rect 20974 35646 21026 35698
rect 22990 35646 23042 35698
rect 23550 35646 23602 35698
rect 25230 35646 25282 35698
rect 27806 35646 27858 35698
rect 28142 35646 28194 35698
rect 28814 35646 28866 35698
rect 34974 35646 35026 35698
rect 37102 35646 37154 35698
rect 38558 35646 38610 35698
rect 39678 35646 39730 35698
rect 3502 35534 3554 35586
rect 6302 35534 6354 35586
rect 8206 35534 8258 35586
rect 10782 35534 10834 35586
rect 11566 35534 11618 35586
rect 13022 35534 13074 35586
rect 14366 35534 14418 35586
rect 15374 35534 15426 35586
rect 23438 35534 23490 35586
rect 25342 35534 25394 35586
rect 26686 35534 26738 35586
rect 27134 35534 27186 35586
rect 29262 35534 29314 35586
rect 41358 35534 41410 35586
rect 12014 35422 12066 35474
rect 4478 35254 4530 35306
rect 4582 35254 4634 35306
rect 4686 35254 4738 35306
rect 35198 35254 35250 35306
rect 35302 35254 35354 35306
rect 35406 35254 35458 35306
rect 12350 35086 12402 35138
rect 2830 34974 2882 35026
rect 9886 34974 9938 35026
rect 17278 34974 17330 35026
rect 18734 34974 18786 35026
rect 20302 34974 20354 35026
rect 26462 34974 26514 35026
rect 26798 34974 26850 35026
rect 27694 34974 27746 35026
rect 29374 34974 29426 35026
rect 30494 34974 30546 35026
rect 6526 34862 6578 34914
rect 8094 34862 8146 34914
rect 8654 34862 8706 34914
rect 10446 34862 10498 34914
rect 10894 34862 10946 34914
rect 12238 34862 12290 34914
rect 12574 34862 12626 34914
rect 13470 34862 13522 34914
rect 14926 34862 14978 34914
rect 16046 34862 16098 34914
rect 16942 34862 16994 34914
rect 19406 34862 19458 34914
rect 20862 34862 20914 34914
rect 22878 34862 22930 34914
rect 23774 34862 23826 34914
rect 25230 34862 25282 34914
rect 26686 34862 26738 34914
rect 27022 34862 27074 34914
rect 27134 34862 27186 34914
rect 27582 34862 27634 34914
rect 27806 34862 27858 34914
rect 29822 34862 29874 34914
rect 30942 34862 30994 34914
rect 32398 34862 32450 34914
rect 32734 34862 32786 34914
rect 35422 34862 35474 34914
rect 36430 34862 36482 34914
rect 38558 34862 38610 34914
rect 39006 34862 39058 34914
rect 2270 34750 2322 34802
rect 2718 34750 2770 34802
rect 2830 34750 2882 34802
rect 5630 34750 5682 34802
rect 7646 34750 7698 34802
rect 11006 34750 11058 34802
rect 11118 34750 11170 34802
rect 11566 34750 11618 34802
rect 14814 34750 14866 34802
rect 15822 34750 15874 34802
rect 16830 34750 16882 34802
rect 18846 34750 18898 34802
rect 21646 34750 21698 34802
rect 24222 34750 24274 34802
rect 25342 34750 25394 34802
rect 26126 34750 26178 34802
rect 33182 34750 33234 34802
rect 34862 34750 34914 34802
rect 36318 34750 36370 34802
rect 37102 34750 37154 34802
rect 39566 34750 39618 34802
rect 1822 34638 1874 34690
rect 2494 34638 2546 34690
rect 6190 34638 6242 34690
rect 12014 34638 12066 34690
rect 12910 34638 12962 34690
rect 13582 34638 13634 34690
rect 13806 34638 13858 34690
rect 19070 34638 19122 34690
rect 19294 34638 19346 34690
rect 20190 34638 20242 34690
rect 20414 34638 20466 34690
rect 22766 34638 22818 34690
rect 28030 34638 28082 34690
rect 28702 34638 28754 34690
rect 32622 34638 32674 34690
rect 35310 34638 35362 34690
rect 37214 34638 37266 34690
rect 19838 34470 19890 34522
rect 19942 34470 19994 34522
rect 20046 34470 20098 34522
rect 50558 34470 50610 34522
rect 50662 34470 50714 34522
rect 50766 34470 50818 34522
rect 1710 34302 1762 34354
rect 3838 34302 3890 34354
rect 5406 34302 5458 34354
rect 6638 34302 6690 34354
rect 7870 34302 7922 34354
rect 11566 34302 11618 34354
rect 13022 34302 13074 34354
rect 13918 34302 13970 34354
rect 15822 34302 15874 34354
rect 18510 34302 18562 34354
rect 21534 34302 21586 34354
rect 23998 34302 24050 34354
rect 24670 34302 24722 34354
rect 29262 34302 29314 34354
rect 29710 34302 29762 34354
rect 30718 34302 30770 34354
rect 2046 34190 2098 34242
rect 10558 34190 10610 34242
rect 14254 34190 14306 34242
rect 14702 34190 14754 34242
rect 15934 34190 15986 34242
rect 17502 34190 17554 34242
rect 18062 34190 18114 34242
rect 19966 34190 20018 34242
rect 21982 34190 22034 34242
rect 23886 34190 23938 34242
rect 28030 34190 28082 34242
rect 28254 34190 28306 34242
rect 35646 34190 35698 34242
rect 8542 34078 8594 34130
rect 9662 34078 9714 34130
rect 10334 34078 10386 34130
rect 10670 34078 10722 34130
rect 12462 34078 12514 34130
rect 12910 34078 12962 34130
rect 14366 34078 14418 34130
rect 15262 34078 15314 34130
rect 16158 34078 16210 34130
rect 16718 34078 16770 34130
rect 17614 34078 17666 34130
rect 18398 34078 18450 34130
rect 18622 34078 18674 34130
rect 19070 34078 19122 34130
rect 19518 34078 19570 34130
rect 20302 34078 20354 34130
rect 20974 34078 21026 34130
rect 21198 34078 21250 34130
rect 22206 34078 22258 34130
rect 22654 34078 22706 34130
rect 23550 34078 23602 34130
rect 23998 34078 24050 34130
rect 25342 34078 25394 34130
rect 25566 34078 25618 34130
rect 26238 34078 26290 34130
rect 28142 34078 28194 34130
rect 33070 34078 33122 34130
rect 36094 34078 36146 34130
rect 36430 34078 36482 34130
rect 39454 34078 39506 34130
rect 2494 33966 2546 34018
rect 3390 33966 3442 34018
rect 5854 33966 5906 34018
rect 7086 33966 7138 34018
rect 7310 33966 7362 34018
rect 8318 33966 8370 34018
rect 10110 33966 10162 34018
rect 11118 33966 11170 34018
rect 12014 33966 12066 34018
rect 27246 33966 27298 34018
rect 28814 33966 28866 34018
rect 30270 33966 30322 34018
rect 34190 33966 34242 34018
rect 36542 33966 36594 34018
rect 38894 33966 38946 34018
rect 8878 33854 8930 33906
rect 17502 33854 17554 33906
rect 26126 33854 26178 33906
rect 27582 33854 27634 33906
rect 4478 33686 4530 33738
rect 4582 33686 4634 33738
rect 4686 33686 4738 33738
rect 35198 33686 35250 33738
rect 35302 33686 35354 33738
rect 35406 33686 35458 33738
rect 14366 33518 14418 33570
rect 14926 33518 14978 33570
rect 16158 33518 16210 33570
rect 16382 33518 16434 33570
rect 18958 33518 19010 33570
rect 32174 33518 32226 33570
rect 7758 33406 7810 33458
rect 9662 33406 9714 33458
rect 14590 33406 14642 33458
rect 15486 33406 15538 33458
rect 17166 33406 17218 33458
rect 20302 33406 20354 33458
rect 23326 33406 23378 33458
rect 26574 33406 26626 33458
rect 27918 33406 27970 33458
rect 2606 33294 2658 33346
rect 3838 33294 3890 33346
rect 4398 33294 4450 33346
rect 4622 33294 4674 33346
rect 5070 33294 5122 33346
rect 5966 33294 6018 33346
rect 9214 33294 9266 33346
rect 17502 33294 17554 33346
rect 18398 33294 18450 33346
rect 19070 33294 19122 33346
rect 23774 33294 23826 33346
rect 25678 33294 25730 33346
rect 27806 33294 27858 33346
rect 28030 33294 28082 33346
rect 30270 33294 30322 33346
rect 30718 33294 30770 33346
rect 33406 33294 33458 33346
rect 35198 33294 35250 33346
rect 36206 33294 36258 33346
rect 37102 33294 37154 33346
rect 39118 33294 39170 33346
rect 41246 33294 41298 33346
rect 1710 33182 1762 33234
rect 3166 33182 3218 33234
rect 3502 33182 3554 33234
rect 4510 33182 4562 33234
rect 7422 33182 7474 33234
rect 8430 33182 8482 33234
rect 17166 33182 17218 33234
rect 18286 33182 18338 33234
rect 25230 33182 25282 33234
rect 26462 33182 26514 33234
rect 28254 33182 28306 33234
rect 29262 33182 29314 33234
rect 32958 33182 33010 33234
rect 33854 33182 33906 33234
rect 38670 33182 38722 33234
rect 40126 33182 40178 33234
rect 2046 33070 2098 33122
rect 3614 33070 3666 33122
rect 10110 33070 10162 33122
rect 12126 33070 12178 33122
rect 12462 33070 12514 33122
rect 13022 33070 13074 33122
rect 13694 33070 13746 33122
rect 14142 33070 14194 33122
rect 15038 33070 15090 33122
rect 16382 33070 16434 33122
rect 18958 33070 19010 33122
rect 19518 33070 19570 33122
rect 20750 33070 20802 33122
rect 21646 33070 21698 33122
rect 22094 33070 22146 33122
rect 22542 33070 22594 33122
rect 22990 33070 23042 33122
rect 23214 33070 23266 33122
rect 23438 33070 23490 33122
rect 27694 33070 27746 33122
rect 36430 33070 36482 33122
rect 37214 33070 37266 33122
rect 37662 33070 37714 33122
rect 19838 32902 19890 32954
rect 19942 32902 19994 32954
rect 20046 32902 20098 32954
rect 50558 32902 50610 32954
rect 50662 32902 50714 32954
rect 50766 32902 50818 32954
rect 6750 32734 6802 32786
rect 13470 32734 13522 32786
rect 19182 32734 19234 32786
rect 28926 32734 28978 32786
rect 34078 32734 34130 32786
rect 40910 32734 40962 32786
rect 5406 32622 5458 32674
rect 13918 32622 13970 32674
rect 14254 32622 14306 32674
rect 18062 32622 18114 32674
rect 21870 32622 21922 32674
rect 22318 32622 22370 32674
rect 22766 32622 22818 32674
rect 28366 32622 28418 32674
rect 28478 32622 28530 32674
rect 33182 32622 33234 32674
rect 35646 32622 35698 32674
rect 37326 32622 37378 32674
rect 41470 32622 41522 32674
rect 2942 32510 2994 32562
rect 3278 32510 3330 32562
rect 3614 32510 3666 32562
rect 4958 32510 5010 32562
rect 6526 32510 6578 32562
rect 7310 32510 7362 32562
rect 8990 32510 9042 32562
rect 10446 32510 10498 32562
rect 12798 32510 12850 32562
rect 13134 32510 13186 32562
rect 16830 32510 16882 32562
rect 17726 32510 17778 32562
rect 18846 32510 18898 32562
rect 21646 32510 21698 32562
rect 23662 32510 23714 32562
rect 25342 32510 25394 32562
rect 27694 32510 27746 32562
rect 28142 32510 28194 32562
rect 34638 32510 34690 32562
rect 35198 32510 35250 32562
rect 38446 32510 38498 32562
rect 38782 32510 38834 32562
rect 8542 32398 8594 32450
rect 10670 32398 10722 32450
rect 14702 32398 14754 32450
rect 15262 32398 15314 32450
rect 16494 32398 16546 32450
rect 18062 32398 18114 32450
rect 19854 32398 19906 32450
rect 21422 32398 21474 32450
rect 24670 32398 24722 32450
rect 27806 32398 27858 32450
rect 39454 32398 39506 32450
rect 10782 32286 10834 32338
rect 26798 32286 26850 32338
rect 4478 32118 4530 32170
rect 4582 32118 4634 32170
rect 4686 32118 4738 32170
rect 35198 32118 35250 32170
rect 35302 32118 35354 32170
rect 35406 32118 35458 32170
rect 17054 31950 17106 32002
rect 25006 31950 25058 32002
rect 2942 31838 2994 31890
rect 3726 31838 3778 31890
rect 15150 31838 15202 31890
rect 20862 31838 20914 31890
rect 23438 31838 23490 31890
rect 27134 31838 27186 31890
rect 29150 31838 29202 31890
rect 30382 31838 30434 31890
rect 33854 31838 33906 31890
rect 3278 31726 3330 31778
rect 4286 31726 4338 31778
rect 8990 31726 9042 31778
rect 9326 31726 9378 31778
rect 9662 31726 9714 31778
rect 11006 31726 11058 31778
rect 12798 31726 12850 31778
rect 13470 31726 13522 31778
rect 14030 31726 14082 31778
rect 14814 31726 14866 31778
rect 15038 31726 15090 31778
rect 15822 31726 15874 31778
rect 16606 31726 16658 31778
rect 17054 31726 17106 31778
rect 17614 31726 17666 31778
rect 18510 31726 18562 31778
rect 19518 31726 19570 31778
rect 20078 31726 20130 31778
rect 20190 31726 20242 31778
rect 20526 31726 20578 31778
rect 22318 31726 22370 31778
rect 22766 31726 22818 31778
rect 25006 31726 25058 31778
rect 26798 31726 26850 31778
rect 28254 31726 28306 31778
rect 33742 31726 33794 31778
rect 34190 31726 34242 31778
rect 38670 31726 38722 31778
rect 39118 31726 39170 31778
rect 11902 31614 11954 31666
rect 14590 31614 14642 31666
rect 16046 31614 16098 31666
rect 17726 31614 17778 31666
rect 21422 31614 21474 31666
rect 24222 31614 24274 31666
rect 25230 31614 25282 31666
rect 27806 31614 27858 31666
rect 28030 31614 28082 31666
rect 33182 31614 33234 31666
rect 35198 31614 35250 31666
rect 36990 31614 37042 31666
rect 39678 31614 39730 31666
rect 12910 31502 12962 31554
rect 15150 31502 15202 31554
rect 18062 31502 18114 31554
rect 18958 31502 19010 31554
rect 19742 31502 19794 31554
rect 20302 31502 20354 31554
rect 29710 31502 29762 31554
rect 30942 31502 30994 31554
rect 37214 31502 37266 31554
rect 19838 31334 19890 31386
rect 19942 31334 19994 31386
rect 20046 31334 20098 31386
rect 50558 31334 50610 31386
rect 50662 31334 50714 31386
rect 50766 31334 50818 31386
rect 2270 31166 2322 31218
rect 7534 31166 7586 31218
rect 9102 31166 9154 31218
rect 10894 31166 10946 31218
rect 13134 31166 13186 31218
rect 14142 31166 14194 31218
rect 15150 31166 15202 31218
rect 16270 31166 16322 31218
rect 17838 31166 17890 31218
rect 18062 31166 18114 31218
rect 18734 31166 18786 31218
rect 19070 31166 19122 31218
rect 20974 31166 21026 31218
rect 23886 31166 23938 31218
rect 25790 31166 25842 31218
rect 26126 31166 26178 31218
rect 26350 31166 26402 31218
rect 26574 31166 26626 31218
rect 27582 31166 27634 31218
rect 27806 31166 27858 31218
rect 27918 31166 27970 31218
rect 28926 31166 28978 31218
rect 33182 31166 33234 31218
rect 3054 31054 3106 31106
rect 4398 31054 4450 31106
rect 5630 31054 5682 31106
rect 12574 31054 12626 31106
rect 13918 31054 13970 31106
rect 15486 31054 15538 31106
rect 17390 31054 17442 31106
rect 17614 31054 17666 31106
rect 18510 31054 18562 31106
rect 18846 31054 18898 31106
rect 20078 31054 20130 31106
rect 20302 31054 20354 31106
rect 21086 31054 21138 31106
rect 21310 31054 21362 31106
rect 24446 31054 24498 31106
rect 24670 31054 24722 31106
rect 34302 31054 34354 31106
rect 35758 31054 35810 31106
rect 2046 30942 2098 30994
rect 3502 30942 3554 30994
rect 4846 30942 4898 30994
rect 5518 30942 5570 30994
rect 10110 30942 10162 30994
rect 11006 30942 11058 30994
rect 11790 30942 11842 30994
rect 13358 30942 13410 30994
rect 14366 30942 14418 30994
rect 14590 30942 14642 30994
rect 16158 30942 16210 30994
rect 16830 30942 16882 30994
rect 18062 30942 18114 30994
rect 18958 30942 19010 30994
rect 20638 30942 20690 30994
rect 24222 30942 24274 30994
rect 26238 30942 26290 30994
rect 28030 30942 28082 30994
rect 28702 30942 28754 30994
rect 29374 30942 29426 30994
rect 34750 30942 34802 30994
rect 36878 30942 36930 30994
rect 38222 30942 38274 30994
rect 3390 30830 3442 30882
rect 6302 30830 6354 30882
rect 8654 30830 8706 30882
rect 14254 30830 14306 30882
rect 19630 30830 19682 30882
rect 21422 30830 21474 30882
rect 21870 30830 21922 30882
rect 24558 30830 24610 30882
rect 25342 30830 25394 30882
rect 27134 30830 27186 30882
rect 8654 30718 8706 30770
rect 9102 30718 9154 30770
rect 16270 30718 16322 30770
rect 27470 30830 27522 30882
rect 28814 30830 28866 30882
rect 37438 30830 37490 30882
rect 20862 30718 20914 30770
rect 21086 30718 21138 30770
rect 21870 30718 21922 30770
rect 27246 30718 27298 30770
rect 4478 30550 4530 30602
rect 4582 30550 4634 30602
rect 4686 30550 4738 30602
rect 35198 30550 35250 30602
rect 35302 30550 35354 30602
rect 35406 30550 35458 30602
rect 4958 30382 5010 30434
rect 14366 30382 14418 30434
rect 14702 30382 14754 30434
rect 21422 30382 21474 30434
rect 6638 30270 6690 30322
rect 11566 30270 11618 30322
rect 14702 30270 14754 30322
rect 15262 30270 15314 30322
rect 17166 30270 17218 30322
rect 26350 30270 26402 30322
rect 27134 30270 27186 30322
rect 28366 30270 28418 30322
rect 30494 30270 30546 30322
rect 31502 30270 31554 30322
rect 34526 30270 34578 30322
rect 1710 30158 1762 30210
rect 6862 30158 6914 30210
rect 7870 30158 7922 30210
rect 8654 30158 8706 30210
rect 9102 30158 9154 30210
rect 9886 30158 9938 30210
rect 11454 30158 11506 30210
rect 12910 30158 12962 30210
rect 17502 30158 17554 30210
rect 17726 30158 17778 30210
rect 20078 30158 20130 30210
rect 21534 30158 21586 30210
rect 21758 30158 21810 30210
rect 22542 30158 22594 30210
rect 23550 30158 23602 30210
rect 25118 30158 25170 30210
rect 25230 30158 25282 30210
rect 25566 30158 25618 30210
rect 30942 30158 30994 30210
rect 31950 30158 32002 30210
rect 34974 30158 35026 30210
rect 35646 30158 35698 30210
rect 37214 30158 37266 30210
rect 2046 30046 2098 30098
rect 2382 30046 2434 30098
rect 5070 30046 5122 30098
rect 6190 30046 6242 30098
rect 6638 30046 6690 30098
rect 7534 30046 7586 30098
rect 9662 30046 9714 30098
rect 11678 30046 11730 30098
rect 12126 30046 12178 30098
rect 12574 30046 12626 30098
rect 19966 30046 20018 30098
rect 21310 30046 21362 30098
rect 21982 30046 22034 30098
rect 22654 30046 22706 30098
rect 23214 30046 23266 30098
rect 24110 30046 24162 30098
rect 24558 30046 24610 30098
rect 25342 30046 25394 30098
rect 35982 30046 36034 30098
rect 36542 30046 36594 30098
rect 2718 29934 2770 29986
rect 3166 29934 3218 29986
rect 4174 29934 4226 29986
rect 4622 29934 4674 29986
rect 4958 29934 5010 29986
rect 5854 29934 5906 29986
rect 6414 29934 6466 29986
rect 7758 29934 7810 29986
rect 10670 29934 10722 29986
rect 11230 29934 11282 29986
rect 11902 29934 11954 29986
rect 12686 29934 12738 29986
rect 13582 29934 13634 29986
rect 14254 29934 14306 29986
rect 19182 29934 19234 29986
rect 23998 29934 24050 29986
rect 26014 29934 26066 29986
rect 29262 29934 29314 29986
rect 19838 29766 19890 29818
rect 19942 29766 19994 29818
rect 20046 29766 20098 29818
rect 50558 29766 50610 29818
rect 50662 29766 50714 29818
rect 50766 29766 50818 29818
rect 1822 29598 1874 29650
rect 6190 29598 6242 29650
rect 7086 29598 7138 29650
rect 15150 29598 15202 29650
rect 18958 29598 19010 29650
rect 19518 29598 19570 29650
rect 20078 29598 20130 29650
rect 23550 29598 23602 29650
rect 23886 29598 23938 29650
rect 24110 29598 24162 29650
rect 24334 29598 24386 29650
rect 25902 29598 25954 29650
rect 27134 29598 27186 29650
rect 27694 29598 27746 29650
rect 35758 29598 35810 29650
rect 3166 29486 3218 29538
rect 6414 29486 6466 29538
rect 7422 29486 7474 29538
rect 9774 29486 9826 29538
rect 11790 29486 11842 29538
rect 13694 29486 13746 29538
rect 13918 29486 13970 29538
rect 14702 29486 14754 29538
rect 20414 29486 20466 29538
rect 22430 29486 22482 29538
rect 29598 29486 29650 29538
rect 34302 29486 34354 29538
rect 37438 29486 37490 29538
rect 2270 29374 2322 29426
rect 4622 29374 4674 29426
rect 5742 29374 5794 29426
rect 7534 29374 7586 29426
rect 7982 29374 8034 29426
rect 8878 29374 8930 29426
rect 9662 29374 9714 29426
rect 10222 29374 10274 29426
rect 11006 29374 11058 29426
rect 12462 29374 12514 29426
rect 13358 29374 13410 29426
rect 14366 29374 14418 29426
rect 14590 29374 14642 29426
rect 19742 29374 19794 29426
rect 19966 29374 20018 29426
rect 20190 29374 20242 29426
rect 20974 29374 21026 29426
rect 21534 29374 21586 29426
rect 21982 29374 22034 29426
rect 24446 29374 24498 29426
rect 27246 29374 27298 29426
rect 27918 29374 27970 29426
rect 28366 29374 28418 29426
rect 28814 29374 28866 29426
rect 29486 29374 29538 29426
rect 35870 29374 35922 29426
rect 38110 29374 38162 29426
rect 12126 29262 12178 29314
rect 15598 29262 15650 29314
rect 26574 29262 26626 29314
rect 27806 29262 27858 29314
rect 10222 29150 10274 29202
rect 13134 29150 13186 29202
rect 13806 29150 13858 29202
rect 29038 29150 29090 29202
rect 4478 28982 4530 29034
rect 4582 28982 4634 29034
rect 4686 28982 4738 29034
rect 35198 28982 35250 29034
rect 35302 28982 35354 29034
rect 35406 28982 35458 29034
rect 21422 28814 21474 28866
rect 30158 28814 30210 28866
rect 2606 28702 2658 28754
rect 3838 28702 3890 28754
rect 10782 28702 10834 28754
rect 11902 28702 11954 28754
rect 12238 28702 12290 28754
rect 12686 28702 12738 28754
rect 15038 28702 15090 28754
rect 16718 28702 16770 28754
rect 18174 28702 18226 28754
rect 19182 28702 19234 28754
rect 20078 28702 20130 28754
rect 26350 28702 26402 28754
rect 26910 28702 26962 28754
rect 27358 28702 27410 28754
rect 2382 28590 2434 28642
rect 2830 28590 2882 28642
rect 3950 28590 4002 28642
rect 6190 28590 6242 28642
rect 6526 28590 6578 28642
rect 10222 28590 10274 28642
rect 11342 28590 11394 28642
rect 14478 28590 14530 28642
rect 15262 28590 15314 28642
rect 15822 28590 15874 28642
rect 16158 28590 16210 28642
rect 18734 28590 18786 28642
rect 20414 28590 20466 28642
rect 20750 28590 20802 28642
rect 21870 28590 21922 28642
rect 22318 28590 22370 28642
rect 22878 28590 22930 28642
rect 23550 28590 23602 28642
rect 24110 28590 24162 28642
rect 25118 28590 25170 28642
rect 26014 28590 26066 28642
rect 28478 28590 28530 28642
rect 29150 28590 29202 28642
rect 29262 28590 29314 28642
rect 29598 28590 29650 28642
rect 29710 28590 29762 28642
rect 3278 28478 3330 28530
rect 7086 28478 7138 28530
rect 10334 28478 10386 28530
rect 11118 28478 11170 28530
rect 14702 28478 14754 28530
rect 14926 28478 14978 28530
rect 18622 28478 18674 28530
rect 21534 28478 21586 28530
rect 23438 28478 23490 28530
rect 24222 28478 24274 28530
rect 28142 28478 28194 28530
rect 28254 28478 28306 28530
rect 2494 28366 2546 28418
rect 2718 28366 2770 28418
rect 3502 28366 3554 28418
rect 3726 28366 3778 28418
rect 4398 28366 4450 28418
rect 7982 28366 8034 28418
rect 10782 28366 10834 28418
rect 10894 28366 10946 28418
rect 15150 28366 15202 28418
rect 18398 28366 18450 28418
rect 20526 28366 20578 28418
rect 21422 28366 21474 28418
rect 24334 28366 24386 28418
rect 27918 28366 27970 28418
rect 19838 28198 19890 28250
rect 19942 28198 19994 28250
rect 20046 28198 20098 28250
rect 50558 28198 50610 28250
rect 50662 28198 50714 28250
rect 50766 28198 50818 28250
rect 2046 28030 2098 28082
rect 3950 28030 4002 28082
rect 4846 28030 4898 28082
rect 5294 28030 5346 28082
rect 7198 28030 7250 28082
rect 8542 28030 8594 28082
rect 8654 28030 8706 28082
rect 8766 28030 8818 28082
rect 11566 28030 11618 28082
rect 13022 28030 13074 28082
rect 18174 28030 18226 28082
rect 18398 28030 18450 28082
rect 25342 28030 25394 28082
rect 25678 28030 25730 28082
rect 27022 28030 27074 28082
rect 29710 28030 29762 28082
rect 30606 28030 30658 28082
rect 3726 27918 3778 27970
rect 5070 27918 5122 27970
rect 6078 27918 6130 27970
rect 7982 27918 8034 27970
rect 8990 27918 9042 27970
rect 12350 27918 12402 27970
rect 16718 27918 16770 27970
rect 20526 27918 20578 27970
rect 20974 27918 21026 27970
rect 21646 27918 21698 27970
rect 27358 27918 27410 27970
rect 1710 27806 1762 27858
rect 4286 27806 4338 27858
rect 5518 27806 5570 27858
rect 5854 27806 5906 27858
rect 6750 27806 6802 27858
rect 7086 27806 7138 27858
rect 7758 27806 7810 27858
rect 8430 27806 8482 27858
rect 10782 27806 10834 27858
rect 12126 27806 12178 27858
rect 13694 27806 13746 27858
rect 14254 27806 14306 27858
rect 15486 27806 15538 27858
rect 15710 27806 15762 27858
rect 15822 27806 15874 27858
rect 16606 27806 16658 27858
rect 17726 27806 17778 27858
rect 17950 27806 18002 27858
rect 18398 27806 18450 27858
rect 18734 27806 18786 27858
rect 19406 27806 19458 27858
rect 19966 27806 20018 27858
rect 20414 27806 20466 27858
rect 25230 27806 25282 27858
rect 25454 27806 25506 27858
rect 26462 27806 26514 27858
rect 26686 27806 26738 27858
rect 27582 27806 27634 27858
rect 30046 27806 30098 27858
rect 2494 27694 2546 27746
rect 3390 27694 3442 27746
rect 3950 27694 4002 27746
rect 5406 27694 5458 27746
rect 9998 27694 10050 27746
rect 22654 27694 22706 27746
rect 24670 27694 24722 27746
rect 28142 27694 28194 27746
rect 29150 27694 29202 27746
rect 16270 27582 16322 27634
rect 16718 27582 16770 27634
rect 19294 27582 19346 27634
rect 4478 27414 4530 27466
rect 4582 27414 4634 27466
rect 4686 27414 4738 27466
rect 35198 27414 35250 27466
rect 35302 27414 35354 27466
rect 35406 27414 35458 27466
rect 15822 27246 15874 27298
rect 24782 27246 24834 27298
rect 6414 27134 6466 27186
rect 8878 27134 8930 27186
rect 9214 27134 9266 27186
rect 10558 27134 10610 27186
rect 12686 27134 12738 27186
rect 14142 27134 14194 27186
rect 14478 27134 14530 27186
rect 17166 27134 17218 27186
rect 17502 27134 17554 27186
rect 17950 27134 18002 27186
rect 18398 27134 18450 27186
rect 19294 27134 19346 27186
rect 20190 27134 20242 27186
rect 23774 27134 23826 27186
rect 26574 27134 26626 27186
rect 27134 27134 27186 27186
rect 5966 27022 6018 27074
rect 9102 27022 9154 27074
rect 9774 27022 9826 27074
rect 12238 27022 12290 27074
rect 13582 27022 13634 27074
rect 14702 27022 14754 27074
rect 15374 27022 15426 27074
rect 15710 27022 15762 27074
rect 18510 27022 18562 27074
rect 18846 27022 18898 27074
rect 24222 27022 24274 27074
rect 24446 27022 24498 27074
rect 25230 27022 25282 27074
rect 26126 27022 26178 27074
rect 4734 26910 4786 26962
rect 10110 26910 10162 26962
rect 15150 26910 15202 26962
rect 15262 26910 15314 26962
rect 18286 26910 18338 26962
rect 25790 26910 25842 26962
rect 9326 26798 9378 26850
rect 15822 26798 15874 26850
rect 16606 26798 16658 26850
rect 21870 26798 21922 26850
rect 19838 26630 19890 26682
rect 19942 26630 19994 26682
rect 20046 26630 20098 26682
rect 50558 26630 50610 26682
rect 50662 26630 50714 26682
rect 50766 26630 50818 26682
rect 6974 26462 7026 26514
rect 7310 26462 7362 26514
rect 9662 26462 9714 26514
rect 9774 26462 9826 26514
rect 10558 26462 10610 26514
rect 12798 26462 12850 26514
rect 13246 26462 13298 26514
rect 13694 26462 13746 26514
rect 14702 26462 14754 26514
rect 15038 26462 15090 26514
rect 15598 26462 15650 26514
rect 15710 26462 15762 26514
rect 17726 26462 17778 26514
rect 25902 26462 25954 26514
rect 26462 26462 26514 26514
rect 7870 26350 7922 26402
rect 11006 26350 11058 26402
rect 15374 26350 15426 26402
rect 17614 26350 17666 26402
rect 18510 26350 18562 26402
rect 5518 26238 5570 26290
rect 5966 26238 6018 26290
rect 9550 26238 9602 26290
rect 10222 26238 10274 26290
rect 11342 26238 11394 26290
rect 11902 26238 11954 26290
rect 12238 26238 12290 26290
rect 15822 26238 15874 26290
rect 16046 26238 16098 26290
rect 17390 26238 17442 26290
rect 17838 26238 17890 26290
rect 17950 26238 18002 26290
rect 21086 26238 21138 26290
rect 21646 26238 21698 26290
rect 22094 26238 22146 26290
rect 14142 26126 14194 26178
rect 16830 26126 16882 26178
rect 19070 26126 19122 26178
rect 19854 26126 19906 26178
rect 20302 26126 20354 26178
rect 20750 26126 20802 26178
rect 22654 26126 22706 26178
rect 23102 26126 23154 26178
rect 25454 26126 25506 26178
rect 4478 25846 4530 25898
rect 4582 25846 4634 25898
rect 4686 25846 4738 25898
rect 35198 25846 35250 25898
rect 35302 25846 35354 25898
rect 35406 25846 35458 25898
rect 7310 25678 7362 25730
rect 7086 25566 7138 25618
rect 8654 25566 8706 25618
rect 13918 25566 13970 25618
rect 16494 25566 16546 25618
rect 17726 25566 17778 25618
rect 18062 25566 18114 25618
rect 19966 25566 20018 25618
rect 23438 25566 23490 25618
rect 27134 25566 27186 25618
rect 28254 25566 28306 25618
rect 7534 25454 7586 25506
rect 7646 25454 7698 25506
rect 8990 25454 9042 25506
rect 9438 25454 9490 25506
rect 9662 25454 9714 25506
rect 10222 25454 10274 25506
rect 10446 25454 10498 25506
rect 11006 25454 11058 25506
rect 11790 25454 11842 25506
rect 11902 25454 11954 25506
rect 12014 25454 12066 25506
rect 12350 25454 12402 25506
rect 12910 25454 12962 25506
rect 14478 25454 14530 25506
rect 15598 25454 15650 25506
rect 16046 25454 16098 25506
rect 17390 25454 17442 25506
rect 18398 25454 18450 25506
rect 18846 25454 18898 25506
rect 19742 25454 19794 25506
rect 20078 25454 20130 25506
rect 21758 25454 21810 25506
rect 23662 25454 23714 25506
rect 25342 25454 25394 25506
rect 25566 25454 25618 25506
rect 1710 25342 1762 25394
rect 2046 25342 2098 25394
rect 2494 25342 2546 25394
rect 7870 25342 7922 25394
rect 9550 25342 9602 25394
rect 10782 25342 10834 25394
rect 12574 25342 12626 25394
rect 14702 25342 14754 25394
rect 16270 25342 16322 25394
rect 20414 25342 20466 25394
rect 22430 25342 22482 25394
rect 23550 25342 23602 25394
rect 9886 25230 9938 25282
rect 11342 25230 11394 25282
rect 12798 25230 12850 25282
rect 13470 25230 13522 25282
rect 15262 25230 15314 25282
rect 18622 25230 18674 25282
rect 21534 25230 21586 25282
rect 27806 25230 27858 25282
rect 29262 25230 29314 25282
rect 19838 25062 19890 25114
rect 19942 25062 19994 25114
rect 20046 25062 20098 25114
rect 50558 25062 50610 25114
rect 50662 25062 50714 25114
rect 50766 25062 50818 25114
rect 6974 24894 7026 24946
rect 7198 24894 7250 24946
rect 8318 24894 8370 24946
rect 11230 24894 11282 24946
rect 11678 24894 11730 24946
rect 16718 24894 16770 24946
rect 17614 24894 17666 24946
rect 22766 24894 22818 24946
rect 25790 24894 25842 24946
rect 26238 24894 26290 24946
rect 16046 24782 16098 24834
rect 19294 24782 19346 24834
rect 20414 24782 20466 24834
rect 22094 24782 22146 24834
rect 24222 24782 24274 24834
rect 7758 24670 7810 24722
rect 12910 24670 12962 24722
rect 13358 24670 13410 24722
rect 13582 24670 13634 24722
rect 13918 24670 13970 24722
rect 16494 24670 16546 24722
rect 17838 24670 17890 24722
rect 21086 24670 21138 24722
rect 22318 24670 22370 24722
rect 24446 24670 24498 24722
rect 18510 24558 18562 24610
rect 25230 24558 25282 24610
rect 4478 24278 4530 24330
rect 4582 24278 4634 24330
rect 4686 24278 4738 24330
rect 35198 24278 35250 24330
rect 35302 24278 35354 24330
rect 35406 24278 35458 24330
rect 20750 24110 20802 24162
rect 11678 23998 11730 24050
rect 13022 23998 13074 24050
rect 14030 23998 14082 24050
rect 15150 23998 15202 24050
rect 16158 23998 16210 24050
rect 19742 23998 19794 24050
rect 21870 23998 21922 24050
rect 23326 23998 23378 24050
rect 24334 23998 24386 24050
rect 25230 23998 25282 24050
rect 25790 23998 25842 24050
rect 14702 23886 14754 23938
rect 15486 23886 15538 23938
rect 16382 23886 16434 23938
rect 18062 23886 18114 23938
rect 19966 23886 20018 23938
rect 20190 23886 20242 23938
rect 20302 23886 20354 23938
rect 21982 23886 22034 23938
rect 22318 23886 22370 23938
rect 23774 23886 23826 23938
rect 24782 23886 24834 23938
rect 1710 23774 1762 23826
rect 2046 23774 2098 23826
rect 16942 23774 16994 23826
rect 18174 23774 18226 23826
rect 21310 23774 21362 23826
rect 2494 23662 2546 23714
rect 19838 23494 19890 23546
rect 19942 23494 19994 23546
rect 20046 23494 20098 23546
rect 50558 23494 50610 23546
rect 50662 23494 50714 23546
rect 50766 23494 50818 23546
rect 15598 23326 15650 23378
rect 15934 23326 15986 23378
rect 16158 23326 16210 23378
rect 16718 23326 16770 23378
rect 18622 23326 18674 23378
rect 19070 23326 19122 23378
rect 21086 23326 21138 23378
rect 21646 23326 21698 23378
rect 22206 23326 22258 23378
rect 22990 23326 23042 23378
rect 25454 23326 25506 23378
rect 15822 23214 15874 23266
rect 19182 23214 19234 23266
rect 21310 23214 21362 23266
rect 15150 22990 15202 23042
rect 17614 22990 17666 23042
rect 19070 22878 19122 22930
rect 4478 22710 4530 22762
rect 4582 22710 4634 22762
rect 4686 22710 4738 22762
rect 35198 22710 35250 22762
rect 35302 22710 35354 22762
rect 35406 22710 35458 22762
rect 15598 22430 15650 22482
rect 1710 22206 1762 22258
rect 2046 22206 2098 22258
rect 2494 22094 2546 22146
rect 19838 21926 19890 21978
rect 19942 21926 19994 21978
rect 20046 21926 20098 21978
rect 50558 21926 50610 21978
rect 50662 21926 50714 21978
rect 50766 21926 50818 21978
rect 4478 21142 4530 21194
rect 4582 21142 4634 21194
rect 4686 21142 4738 21194
rect 35198 21142 35250 21194
rect 35302 21142 35354 21194
rect 35406 21142 35458 21194
rect 2046 20638 2098 20690
rect 1710 20526 1762 20578
rect 2494 20526 2546 20578
rect 19838 20358 19890 20410
rect 19942 20358 19994 20410
rect 20046 20358 20098 20410
rect 50558 20358 50610 20410
rect 50662 20358 50714 20410
rect 50766 20358 50818 20410
rect 4478 19574 4530 19626
rect 4582 19574 4634 19626
rect 4686 19574 4738 19626
rect 35198 19574 35250 19626
rect 35302 19574 35354 19626
rect 35406 19574 35458 19626
rect 19838 18790 19890 18842
rect 19942 18790 19994 18842
rect 20046 18790 20098 18842
rect 50558 18790 50610 18842
rect 50662 18790 50714 18842
rect 50766 18790 50818 18842
rect 2046 18622 2098 18674
rect 1710 18398 1762 18450
rect 2494 18286 2546 18338
rect 4478 18006 4530 18058
rect 4582 18006 4634 18058
rect 4686 18006 4738 18058
rect 35198 18006 35250 18058
rect 35302 18006 35354 18058
rect 35406 18006 35458 18058
rect 19838 17222 19890 17274
rect 19942 17222 19994 17274
rect 20046 17222 20098 17274
rect 50558 17222 50610 17274
rect 50662 17222 50714 17274
rect 50766 17222 50818 17274
rect 2046 17054 2098 17106
rect 1710 16830 1762 16882
rect 2494 16830 2546 16882
rect 4478 16438 4530 16490
rect 4582 16438 4634 16490
rect 4686 16438 4738 16490
rect 35198 16438 35250 16490
rect 35302 16438 35354 16490
rect 35406 16438 35458 16490
rect 19838 15654 19890 15706
rect 19942 15654 19994 15706
rect 20046 15654 20098 15706
rect 50558 15654 50610 15706
rect 50662 15654 50714 15706
rect 50766 15654 50818 15706
rect 2046 15486 2098 15538
rect 1710 15262 1762 15314
rect 2494 15150 2546 15202
rect 4478 14870 4530 14922
rect 4582 14870 4634 14922
rect 4686 14870 4738 14922
rect 35198 14870 35250 14922
rect 35302 14870 35354 14922
rect 35406 14870 35458 14922
rect 19838 14086 19890 14138
rect 19942 14086 19994 14138
rect 20046 14086 20098 14138
rect 50558 14086 50610 14138
rect 50662 14086 50714 14138
rect 50766 14086 50818 14138
rect 4478 13302 4530 13354
rect 4582 13302 4634 13354
rect 4686 13302 4738 13354
rect 35198 13302 35250 13354
rect 35302 13302 35354 13354
rect 35406 13302 35458 13354
rect 1710 12798 1762 12850
rect 2046 12798 2098 12850
rect 2494 12798 2546 12850
rect 19838 12518 19890 12570
rect 19942 12518 19994 12570
rect 20046 12518 20098 12570
rect 50558 12518 50610 12570
rect 50662 12518 50714 12570
rect 50766 12518 50818 12570
rect 4478 11734 4530 11786
rect 4582 11734 4634 11786
rect 4686 11734 4738 11786
rect 35198 11734 35250 11786
rect 35302 11734 35354 11786
rect 35406 11734 35458 11786
rect 1710 11230 1762 11282
rect 2046 11230 2098 11282
rect 2494 11118 2546 11170
rect 19838 10950 19890 11002
rect 19942 10950 19994 11002
rect 20046 10950 20098 11002
rect 50558 10950 50610 11002
rect 50662 10950 50714 11002
rect 50766 10950 50818 11002
rect 4478 10166 4530 10218
rect 4582 10166 4634 10218
rect 4686 10166 4738 10218
rect 35198 10166 35250 10218
rect 35302 10166 35354 10218
rect 35406 10166 35458 10218
rect 1710 9662 1762 9714
rect 2046 9662 2098 9714
rect 2494 9550 2546 9602
rect 19838 9382 19890 9434
rect 19942 9382 19994 9434
rect 20046 9382 20098 9434
rect 50558 9382 50610 9434
rect 50662 9382 50714 9434
rect 50766 9382 50818 9434
rect 4478 8598 4530 8650
rect 4582 8598 4634 8650
rect 4686 8598 4738 8650
rect 35198 8598 35250 8650
rect 35302 8598 35354 8650
rect 35406 8598 35458 8650
rect 1710 8094 1762 8146
rect 2046 8094 2098 8146
rect 2494 7982 2546 8034
rect 19838 7814 19890 7866
rect 19942 7814 19994 7866
rect 20046 7814 20098 7866
rect 50558 7814 50610 7866
rect 50662 7814 50714 7866
rect 50766 7814 50818 7866
rect 4478 7030 4530 7082
rect 4582 7030 4634 7082
rect 4686 7030 4738 7082
rect 35198 7030 35250 7082
rect 35302 7030 35354 7082
rect 35406 7030 35458 7082
rect 19838 6246 19890 6298
rect 19942 6246 19994 6298
rect 20046 6246 20098 6298
rect 50558 6246 50610 6298
rect 50662 6246 50714 6298
rect 50766 6246 50818 6298
rect 1710 5854 1762 5906
rect 2158 5742 2210 5794
rect 4478 5462 4530 5514
rect 4582 5462 4634 5514
rect 4686 5462 4738 5514
rect 35198 5462 35250 5514
rect 35302 5462 35354 5514
rect 35406 5462 35458 5514
rect 1822 5182 1874 5234
rect 19838 4678 19890 4730
rect 19942 4678 19994 4730
rect 20046 4678 20098 4730
rect 50558 4678 50610 4730
rect 50662 4678 50714 4730
rect 50766 4678 50818 4730
rect 2046 4510 2098 4562
rect 1710 4286 1762 4338
rect 2494 4174 2546 4226
rect 4478 3894 4530 3946
rect 4582 3894 4634 3946
rect 4686 3894 4738 3946
rect 35198 3894 35250 3946
rect 35302 3894 35354 3946
rect 35406 3894 35458 3946
rect 2270 3614 2322 3666
rect 1710 3390 1762 3442
rect 2718 3390 2770 3442
rect 19838 3110 19890 3162
rect 19942 3110 19994 3162
rect 20046 3110 20098 3162
rect 50558 3110 50610 3162
rect 50662 3110 50714 3162
rect 50766 3110 50818 3162
<< metal2 >>
rect 2912 59200 3024 60000
rect 5152 59200 5264 60000
rect 7392 59200 7504 60000
rect 9632 59200 9744 60000
rect 11872 59200 11984 60000
rect 14112 59200 14224 60000
rect 16352 59200 16464 60000
rect 18592 59200 18704 60000
rect 20832 59200 20944 60000
rect 23072 59200 23184 60000
rect 25312 59200 25424 60000
rect 27552 59200 27664 60000
rect 29792 59200 29904 60000
rect 32032 59200 32144 60000
rect 34272 59200 34384 60000
rect 36512 59200 36624 60000
rect 38752 59200 38864 60000
rect 40992 59200 41104 60000
rect 43232 59200 43344 60000
rect 45472 59200 45584 60000
rect 47712 59200 47824 60000
rect 49952 59200 50064 60000
rect 52192 59200 52304 60000
rect 54432 59200 54544 60000
rect 56672 59200 56784 60000
rect 2156 57652 2212 57662
rect 2044 56194 2100 56206
rect 2044 56142 2046 56194
rect 2098 56142 2100 56194
rect 1708 56082 1764 56094
rect 1708 56030 1710 56082
rect 1762 56030 1764 56082
rect 1708 55860 1764 56030
rect 1708 55794 1764 55804
rect 2044 55468 2100 56142
rect 1932 55412 2100 55468
rect 2156 56084 2212 57596
rect 1372 54628 1428 54638
rect 1148 39620 1204 39630
rect 1036 35812 1092 35822
rect 1036 23492 1092 35756
rect 1148 29764 1204 39564
rect 1372 36372 1428 54572
rect 1708 54514 1764 54526
rect 1708 54462 1710 54514
rect 1762 54462 1764 54514
rect 1708 54068 1764 54462
rect 1708 54002 1764 54012
rect 1708 52946 1764 52958
rect 1708 52894 1710 52946
rect 1762 52894 1764 52946
rect 1708 52836 1764 52894
rect 1708 52276 1764 52780
rect 1708 52210 1764 52220
rect 1820 51378 1876 51390
rect 1820 51326 1822 51378
rect 1874 51326 1876 51378
rect 1820 51268 1876 51326
rect 1708 50708 1764 50718
rect 1708 50614 1764 50652
rect 1708 50484 1764 50494
rect 1820 50484 1876 51212
rect 1764 50428 1876 50484
rect 1708 50418 1764 50428
rect 1932 49812 1988 55412
rect 2156 55410 2212 56028
rect 2380 56194 2436 56206
rect 2380 56142 2382 56194
rect 2434 56142 2436 56194
rect 2380 55468 2436 56142
rect 2604 56084 2660 56094
rect 2604 55990 2660 56028
rect 2380 55412 2660 55468
rect 2156 55358 2158 55410
rect 2210 55358 2212 55410
rect 2156 55346 2212 55358
rect 2044 54628 2100 54638
rect 2044 54534 2100 54572
rect 2492 54402 2548 54414
rect 2492 54350 2494 54402
rect 2546 54350 2548 54402
rect 2492 54068 2548 54350
rect 2492 54002 2548 54012
rect 2044 53060 2100 53070
rect 2044 53058 2324 53060
rect 2044 53006 2046 53058
rect 2098 53006 2324 53058
rect 2044 53004 2324 53006
rect 2044 52994 2100 53004
rect 2044 51492 2100 51502
rect 2044 51398 2100 51436
rect 2268 50428 2324 53004
rect 2492 52836 2548 52846
rect 2492 52742 2548 52780
rect 2492 51268 2548 51278
rect 2492 51174 2548 51212
rect 2268 50372 2436 50428
rect 1932 49756 2324 49812
rect 1708 49700 1764 49710
rect 1708 49698 2212 49700
rect 1708 49646 1710 49698
rect 1762 49646 2212 49698
rect 1708 49644 2212 49646
rect 1708 49634 1764 49644
rect 1708 48914 1764 48926
rect 1708 48862 1710 48914
rect 1762 48862 1764 48914
rect 1708 48692 1764 48862
rect 2044 48804 2100 48814
rect 1708 48626 1764 48636
rect 1820 48802 2100 48804
rect 1820 48750 2046 48802
rect 2098 48750 2100 48802
rect 1820 48748 2100 48750
rect 1708 46900 1764 46910
rect 1708 46786 1764 46844
rect 1708 46734 1710 46786
rect 1762 46734 1764 46786
rect 1708 46722 1764 46734
rect 1708 45778 1764 45790
rect 1708 45726 1710 45778
rect 1762 45726 1764 45778
rect 1708 45108 1764 45726
rect 1708 45042 1764 45052
rect 1372 36306 1428 36316
rect 1484 44884 1540 44894
rect 1148 29698 1204 29708
rect 1260 32452 1316 32462
rect 1036 23426 1092 23436
rect 1148 26964 1204 26974
rect 1148 15204 1204 26908
rect 1148 15138 1204 15148
rect 1260 5908 1316 32396
rect 1484 28308 1540 44828
rect 1820 43652 1876 48748
rect 2044 48738 2100 48748
rect 2156 47684 2212 49644
rect 2156 47458 2212 47628
rect 2156 47406 2158 47458
rect 2210 47406 2212 47458
rect 2156 47394 2212 47406
rect 2268 47236 2324 49756
rect 2156 47180 2324 47236
rect 2380 47236 2436 50372
rect 2492 48802 2548 48814
rect 2492 48750 2494 48802
rect 2546 48750 2548 48802
rect 2492 48692 2548 48750
rect 2492 48626 2548 48636
rect 2604 47796 2660 55412
rect 2940 53844 2996 59200
rect 5068 56308 5124 56318
rect 5180 56308 5236 59200
rect 7420 56308 7476 59200
rect 7644 56308 7700 56318
rect 5068 56306 5572 56308
rect 5068 56254 5070 56306
rect 5122 56254 5572 56306
rect 5068 56252 5572 56254
rect 5068 56242 5124 56252
rect 5516 56194 5572 56252
rect 7420 56306 7700 56308
rect 7420 56254 7422 56306
rect 7474 56254 7646 56306
rect 7698 56254 7700 56306
rect 7420 56252 7700 56254
rect 7420 56242 7476 56252
rect 7644 56242 7700 56252
rect 9660 56308 9716 59200
rect 9884 56308 9940 56318
rect 9660 56306 9940 56308
rect 9660 56254 9662 56306
rect 9714 56254 9886 56306
rect 9938 56254 9940 56306
rect 9660 56252 9940 56254
rect 9660 56242 9716 56252
rect 9884 56242 9940 56252
rect 11900 56308 11956 59200
rect 14140 56420 14196 59200
rect 14140 56364 14644 56420
rect 12124 56308 12180 56318
rect 11900 56306 12180 56308
rect 11900 56254 11902 56306
rect 11954 56254 12126 56306
rect 12178 56254 12180 56306
rect 11900 56252 12180 56254
rect 11900 56242 11956 56252
rect 12124 56242 12180 56252
rect 14140 56306 14196 56364
rect 14140 56254 14142 56306
rect 14194 56254 14196 56306
rect 14140 56242 14196 56254
rect 5516 56142 5518 56194
rect 5570 56142 5572 56194
rect 5516 56130 5572 56142
rect 5852 56194 5908 56206
rect 5852 56142 5854 56194
rect 5906 56142 5908 56194
rect 3164 55970 3220 55982
rect 3164 55918 3166 55970
rect 3218 55918 3220 55970
rect 3164 55860 3220 55918
rect 3164 55794 3220 55804
rect 4476 55692 4740 55702
rect 4532 55636 4580 55692
rect 4636 55636 4684 55692
rect 4476 55626 4740 55636
rect 5852 55188 5908 56142
rect 7980 56194 8036 56206
rect 7980 56142 7982 56194
rect 8034 56142 8036 56194
rect 7980 55468 8036 56142
rect 10220 56194 10276 56206
rect 10220 56142 10222 56194
rect 10274 56142 10276 56194
rect 10220 55468 10276 56142
rect 12460 56194 12516 56206
rect 12460 56142 12462 56194
rect 12514 56142 12516 56194
rect 12460 55468 12516 56142
rect 14364 56194 14420 56206
rect 14364 56142 14366 56194
rect 14418 56142 14420 56194
rect 14364 55468 14420 56142
rect 14588 56082 14644 56364
rect 16380 56308 16436 59200
rect 16492 56308 16548 56318
rect 16940 56308 16996 56318
rect 16380 56306 16996 56308
rect 16380 56254 16494 56306
rect 16546 56254 16942 56306
rect 16994 56254 16996 56306
rect 16380 56252 16996 56254
rect 16492 56242 16548 56252
rect 16940 56242 16996 56252
rect 18620 56308 18676 59200
rect 19836 56476 20100 56486
rect 19892 56420 19940 56476
rect 19996 56420 20044 56476
rect 19836 56410 20100 56420
rect 18844 56308 18900 56318
rect 18620 56306 18900 56308
rect 18620 56254 18622 56306
rect 18674 56254 18846 56306
rect 18898 56254 18900 56306
rect 18620 56252 18900 56254
rect 18620 56242 18676 56252
rect 18844 56242 18900 56252
rect 20300 56308 20356 56318
rect 20860 56308 20916 59200
rect 20300 56306 20916 56308
rect 20300 56254 20302 56306
rect 20354 56254 20916 56306
rect 20300 56252 20916 56254
rect 20300 56242 20356 56252
rect 17276 56196 17332 56206
rect 17276 56194 17556 56196
rect 17276 56142 17278 56194
rect 17330 56142 17556 56194
rect 17276 56140 17556 56142
rect 17276 56130 17332 56140
rect 14588 56030 14590 56082
rect 14642 56030 14644 56082
rect 14588 56018 14644 56030
rect 7980 55412 8260 55468
rect 10220 55412 10500 55468
rect 12460 55412 12740 55468
rect 5852 55122 5908 55132
rect 4476 54124 4740 54134
rect 4532 54068 4580 54124
rect 4636 54068 4684 54124
rect 4476 54058 4740 54068
rect 2940 53778 2996 53788
rect 5740 53844 5796 53854
rect 4476 52556 4740 52566
rect 4532 52500 4580 52556
rect 4636 52500 4684 52556
rect 4476 52490 4740 52500
rect 3836 51940 3892 51950
rect 2716 51492 2772 51502
rect 2716 50428 2772 51436
rect 3276 50708 3332 50718
rect 2716 50372 2884 50428
rect 2604 47740 2772 47796
rect 2604 47572 2660 47582
rect 2492 47570 2660 47572
rect 2492 47518 2606 47570
rect 2658 47518 2660 47570
rect 2492 47516 2660 47518
rect 2492 47460 2548 47516
rect 2604 47506 2660 47516
rect 2492 47394 2548 47404
rect 2380 47180 2660 47236
rect 2044 46788 2100 46798
rect 1708 43596 1876 43652
rect 1932 46786 2100 46788
rect 1932 46734 2046 46786
rect 2098 46734 2100 46786
rect 1932 46732 2100 46734
rect 1708 42308 1764 43596
rect 1820 43426 1876 43438
rect 1820 43374 1822 43426
rect 1874 43374 1876 43426
rect 1820 43316 1876 43374
rect 1820 42754 1876 43260
rect 1820 42702 1822 42754
rect 1874 42702 1876 42754
rect 1820 42690 1876 42702
rect 1932 42420 1988 46732
rect 2044 46722 2100 46732
rect 2044 45666 2100 45678
rect 2044 45614 2046 45666
rect 2098 45614 2100 45666
rect 2044 43652 2100 45614
rect 2044 43586 2100 43596
rect 2044 43428 2100 43438
rect 2044 42642 2100 43372
rect 2156 43092 2212 47180
rect 2492 46900 2548 46910
rect 2492 46806 2548 46844
rect 2492 45668 2548 45678
rect 2380 45666 2548 45668
rect 2380 45614 2494 45666
rect 2546 45614 2548 45666
rect 2380 45612 2548 45614
rect 2268 45108 2324 45118
rect 2380 45108 2436 45612
rect 2492 45602 2548 45612
rect 2604 45330 2660 47180
rect 2604 45278 2606 45330
rect 2658 45278 2660 45330
rect 2604 45266 2660 45278
rect 2324 45052 2436 45108
rect 2492 45108 2548 45118
rect 2268 45042 2324 45052
rect 2492 44212 2548 45052
rect 2380 44156 2548 44212
rect 2268 44100 2324 44110
rect 2268 43650 2324 44044
rect 2380 43876 2436 44156
rect 2716 44100 2772 47740
rect 2828 46228 2884 50372
rect 3276 48468 3332 50652
rect 3836 50706 3892 51884
rect 4396 51380 4452 51390
rect 4396 51286 4452 51324
rect 5180 51380 5236 51390
rect 5068 51268 5124 51278
rect 5068 51174 5124 51212
rect 4476 50988 4740 50998
rect 4532 50932 4580 50988
rect 4636 50932 4684 50988
rect 4476 50922 4740 50932
rect 5068 50708 5124 50718
rect 5180 50708 5236 51324
rect 3836 50654 3838 50706
rect 3890 50654 3892 50706
rect 3836 50642 3892 50654
rect 4620 50706 5236 50708
rect 4620 50654 5070 50706
rect 5122 50654 5236 50706
rect 4620 50652 5236 50654
rect 4620 50594 4676 50652
rect 4620 50542 4622 50594
rect 4674 50542 4676 50594
rect 3836 49924 3892 49934
rect 3836 49830 3892 49868
rect 4620 49810 4676 50542
rect 5068 50034 5124 50652
rect 5068 49982 5070 50034
rect 5122 49982 5124 50034
rect 5068 49970 5124 49982
rect 4620 49758 4622 49810
rect 4674 49758 4676 49810
rect 4620 49746 4676 49758
rect 4476 49420 4740 49430
rect 4532 49364 4580 49420
rect 4636 49364 4684 49420
rect 4476 49354 4740 49364
rect 3500 48468 3556 48478
rect 3276 48466 3556 48468
rect 3276 48414 3502 48466
rect 3554 48414 3556 48466
rect 3276 48412 3556 48414
rect 3276 47684 3332 47694
rect 3276 47590 3332 47628
rect 3388 47460 3444 48412
rect 3500 48402 3556 48412
rect 4060 48130 4116 48142
rect 4060 48078 4062 48130
rect 4114 48078 4116 48130
rect 3164 47404 3444 47460
rect 3948 47460 4004 47470
rect 3052 47348 3108 47358
rect 3164 47348 3220 47404
rect 2940 47346 3220 47348
rect 2940 47294 3054 47346
rect 3106 47294 3220 47346
rect 2940 47292 3220 47294
rect 2940 46786 2996 47292
rect 3052 47282 3108 47292
rect 2940 46734 2942 46786
rect 2994 46734 2996 46786
rect 2940 46722 2996 46734
rect 3612 47234 3668 47246
rect 3612 47182 3614 47234
rect 3666 47182 3668 47234
rect 3052 46452 3108 46462
rect 3052 46450 3332 46452
rect 3052 46398 3054 46450
rect 3106 46398 3332 46450
rect 3052 46396 3332 46398
rect 3052 46386 3108 46396
rect 2828 46172 3220 46228
rect 3164 45330 3220 46172
rect 3164 45278 3166 45330
rect 3218 45278 3220 45330
rect 3164 45266 3220 45278
rect 2828 45108 2884 45118
rect 3052 45108 3108 45118
rect 2828 45106 2996 45108
rect 2828 45054 2830 45106
rect 2882 45054 2996 45106
rect 2828 45052 2996 45054
rect 2828 45042 2884 45052
rect 2716 44034 2772 44044
rect 2380 43820 2548 43876
rect 2268 43598 2270 43650
rect 2322 43598 2324 43650
rect 2268 43586 2324 43598
rect 2380 43540 2436 43550
rect 2156 43036 2324 43092
rect 2044 42590 2046 42642
rect 2098 42590 2100 42642
rect 2044 42578 2100 42590
rect 1932 42364 2212 42420
rect 1708 42252 1988 42308
rect 1820 41860 1876 41870
rect 1708 41858 1876 41860
rect 1708 41806 1822 41858
rect 1874 41806 1876 41858
rect 1708 41804 1876 41806
rect 1708 41524 1764 41804
rect 1820 41794 1876 41804
rect 1708 41186 1764 41468
rect 1708 41134 1710 41186
rect 1762 41134 1764 41186
rect 1708 41122 1764 41134
rect 1708 40402 1764 40414
rect 1708 40350 1710 40402
rect 1762 40350 1764 40402
rect 1708 40292 1764 40350
rect 1708 39732 1764 40236
rect 1708 39666 1764 39676
rect 1820 38722 1876 38734
rect 1820 38670 1822 38722
rect 1874 38670 1876 38722
rect 1820 38668 1876 38670
rect 1708 38612 1876 38668
rect 1708 37940 1764 38612
rect 1708 37846 1764 37884
rect 1932 37492 1988 42252
rect 2044 41972 2100 41982
rect 2044 41074 2100 41916
rect 2044 41022 2046 41074
rect 2098 41022 2100 41074
rect 2044 41010 2100 41022
rect 2044 40514 2100 40526
rect 2044 40462 2046 40514
rect 2098 40462 2100 40514
rect 2044 39620 2100 40462
rect 2044 39554 2100 39564
rect 2044 37826 2100 37838
rect 2044 37774 2046 37826
rect 2098 37774 2100 37826
rect 2044 37604 2100 37774
rect 2156 37716 2212 42364
rect 2268 42082 2324 43036
rect 2268 42030 2270 42082
rect 2322 42030 2324 42082
rect 2268 42018 2324 42030
rect 2380 41300 2436 43484
rect 2268 41244 2436 41300
rect 2492 43538 2548 43820
rect 2940 43708 2996 45052
rect 3052 45014 3108 45052
rect 3164 44884 3220 44894
rect 3164 44790 3220 44828
rect 3276 43708 3332 46396
rect 2716 43652 2772 43662
rect 2940 43652 3220 43708
rect 3276 43652 3556 43708
rect 2716 43558 2772 43596
rect 2492 43486 2494 43538
rect 2546 43486 2548 43538
rect 2492 41970 2548 43486
rect 2940 43538 2996 43550
rect 2940 43486 2942 43538
rect 2994 43486 2996 43538
rect 2828 43426 2884 43438
rect 2828 43374 2830 43426
rect 2882 43374 2884 43426
rect 2716 42642 2772 42654
rect 2716 42590 2718 42642
rect 2770 42590 2772 42642
rect 2716 42308 2772 42590
rect 2828 42642 2884 43374
rect 2828 42590 2830 42642
rect 2882 42590 2884 42642
rect 2828 42578 2884 42590
rect 2716 42242 2772 42252
rect 2492 41918 2494 41970
rect 2546 41918 2548 41970
rect 2268 39172 2324 41244
rect 2380 41074 2436 41086
rect 2380 41022 2382 41074
rect 2434 41022 2436 41074
rect 2380 39620 2436 41022
rect 2492 41076 2548 41918
rect 2716 41972 2772 41982
rect 2716 41878 2772 41916
rect 2828 41972 2884 41982
rect 2940 41972 2996 43486
rect 3052 42532 3108 42542
rect 3052 42438 3108 42476
rect 2828 41970 2996 41972
rect 2828 41918 2830 41970
rect 2882 41918 2996 41970
rect 2828 41916 2996 41918
rect 3052 42308 3108 42318
rect 2604 41858 2660 41870
rect 2604 41806 2606 41858
rect 2658 41806 2660 41858
rect 2604 41188 2660 41806
rect 2604 41122 2660 41132
rect 2492 41010 2548 41020
rect 2716 41076 2772 41086
rect 2716 40982 2772 41020
rect 2828 40516 2884 41916
rect 3052 40628 3108 42252
rect 3164 40740 3220 43652
rect 3500 43538 3556 43652
rect 3612 43652 3668 47182
rect 3724 47124 3780 47134
rect 3724 46786 3780 47068
rect 3724 46734 3726 46786
rect 3778 46734 3780 46786
rect 3724 46722 3780 46734
rect 3948 46676 4004 47404
rect 4060 47124 4116 48078
rect 4476 47852 4740 47862
rect 4532 47796 4580 47852
rect 4636 47796 4684 47852
rect 4476 47786 4740 47796
rect 4060 47058 4116 47068
rect 4508 47346 4564 47358
rect 4508 47294 4510 47346
rect 4562 47294 4564 47346
rect 4508 46900 4564 47294
rect 5740 47236 5796 53788
rect 7980 52948 8036 52958
rect 7980 52854 8036 52892
rect 5852 52834 5908 52846
rect 5852 52782 5854 52834
rect 5906 52782 5908 52834
rect 5852 50820 5908 52782
rect 7644 51380 7700 51390
rect 7644 51286 7700 51324
rect 7196 51268 7252 51278
rect 5852 50754 5908 50764
rect 7084 51266 7252 51268
rect 7084 51214 7198 51266
rect 7250 51214 7252 51266
rect 7084 51212 7252 51214
rect 7084 50708 7140 51212
rect 7196 51202 7252 51212
rect 7308 50820 7364 50830
rect 6748 50706 7140 50708
rect 6748 50654 7086 50706
rect 7138 50654 7140 50706
rect 6748 50652 7140 50654
rect 6748 50428 6804 50652
rect 7084 50642 7140 50652
rect 7196 50764 7308 50820
rect 6636 50372 6804 50428
rect 6524 49812 6580 49822
rect 6636 49812 6692 50372
rect 6524 49810 6692 49812
rect 6524 49758 6526 49810
rect 6578 49758 6692 49810
rect 6524 49756 6692 49758
rect 6524 49746 6580 49756
rect 6412 49586 6468 49598
rect 6412 49534 6414 49586
rect 6466 49534 6468 49586
rect 5740 47170 5796 47180
rect 6076 48244 6132 48254
rect 6076 48130 6132 48188
rect 6076 48078 6078 48130
rect 6130 48078 6132 48130
rect 4508 46834 4564 46844
rect 4844 46788 4900 46798
rect 4844 46694 4900 46732
rect 4508 46676 4564 46686
rect 3948 46674 4564 46676
rect 3948 46622 3950 46674
rect 4002 46622 4510 46674
rect 4562 46622 4564 46674
rect 3948 46620 4564 46622
rect 3836 46562 3892 46574
rect 3836 46510 3838 46562
rect 3890 46510 3892 46562
rect 3836 45556 3892 46510
rect 3948 45890 4004 46620
rect 4508 46610 4564 46620
rect 5964 46562 6020 46574
rect 5964 46510 5966 46562
rect 6018 46510 6020 46562
rect 4476 46284 4740 46294
rect 4532 46228 4580 46284
rect 4636 46228 4684 46284
rect 4476 46218 4740 46228
rect 3948 45838 3950 45890
rect 4002 45838 4004 45890
rect 3948 45826 4004 45838
rect 4508 45780 4564 45790
rect 4508 45686 4564 45724
rect 3836 45500 4228 45556
rect 4172 45444 4228 45500
rect 4060 45332 4116 45342
rect 3836 45276 4060 45332
rect 3836 44994 3892 45276
rect 3836 44942 3838 44994
rect 3890 44942 3892 44994
rect 3836 44930 3892 44942
rect 3612 43586 3668 43596
rect 3500 43486 3502 43538
rect 3554 43486 3556 43538
rect 3500 42194 3556 43486
rect 3724 43316 3780 43326
rect 3500 42142 3502 42194
rect 3554 42142 3556 42194
rect 3500 42130 3556 42142
rect 3612 43260 3724 43316
rect 3164 40684 3332 40740
rect 3052 40572 3220 40628
rect 2716 40460 2884 40516
rect 2492 40402 2548 40414
rect 2492 40350 2494 40402
rect 2546 40350 2548 40402
rect 2492 40292 2548 40350
rect 2492 40226 2548 40236
rect 2604 39620 2660 39630
rect 2380 39564 2604 39620
rect 2268 39116 2548 39172
rect 2380 38946 2436 38958
rect 2380 38894 2382 38946
rect 2434 38894 2436 38946
rect 2380 38052 2436 38894
rect 2492 38668 2548 39116
rect 2604 38834 2660 39564
rect 2604 38782 2606 38834
rect 2658 38782 2660 38834
rect 2604 38770 2660 38782
rect 2492 38612 2660 38668
rect 2492 38052 2548 38062
rect 2380 38050 2548 38052
rect 2380 37998 2494 38050
rect 2546 37998 2548 38050
rect 2380 37996 2548 37998
rect 2156 37660 2324 37716
rect 2044 37548 2212 37604
rect 1932 37426 1988 37436
rect 2044 37378 2100 37390
rect 2044 37326 2046 37378
rect 2098 37326 2100 37378
rect 1708 37266 1764 37278
rect 1708 37214 1710 37266
rect 1762 37214 1764 37266
rect 1708 37156 1764 37214
rect 1708 36148 1764 37100
rect 2044 36708 2100 37326
rect 1932 36652 2100 36708
rect 1932 36596 1988 36652
rect 1820 36540 1988 36596
rect 1820 36148 1876 36540
rect 2044 36484 2100 36494
rect 1932 36372 1988 36382
rect 1932 36278 1988 36316
rect 1820 36092 1988 36148
rect 1708 36082 1764 36092
rect 1820 34690 1876 34702
rect 1820 34638 1822 34690
rect 1874 34638 1876 34690
rect 1708 34356 1764 34366
rect 1820 34356 1876 34638
rect 1764 34300 1876 34356
rect 1708 34262 1764 34300
rect 1708 33236 1764 33246
rect 1708 32564 1764 33180
rect 1708 32498 1764 32508
rect 1932 31220 1988 36092
rect 2044 34468 2100 36428
rect 2156 34916 2212 37548
rect 2268 35810 2324 37660
rect 2492 37378 2548 37996
rect 2604 37938 2660 38612
rect 2716 38052 2772 40460
rect 2828 40292 2884 40302
rect 2828 39506 2884 40236
rect 2828 39454 2830 39506
rect 2882 39454 2884 39506
rect 2828 39442 2884 39454
rect 3052 39508 3108 39518
rect 3052 39414 3108 39452
rect 2940 39394 2996 39406
rect 2940 39342 2942 39394
rect 2994 39342 2996 39394
rect 2940 38388 2996 39342
rect 2940 38322 2996 38332
rect 3052 38052 3108 38062
rect 2716 38050 3108 38052
rect 2716 37998 3054 38050
rect 3106 37998 3108 38050
rect 2716 37996 3108 37998
rect 2604 37886 2606 37938
rect 2658 37886 2660 37938
rect 2604 37874 2660 37886
rect 2828 37828 2884 37838
rect 2716 37826 2884 37828
rect 2716 37774 2830 37826
rect 2882 37774 2884 37826
rect 2716 37772 2884 37774
rect 2604 37492 2660 37502
rect 2604 37398 2660 37436
rect 2492 37326 2494 37378
rect 2546 37326 2548 37378
rect 2492 36482 2548 37326
rect 2716 36708 2772 37772
rect 2828 37762 2884 37772
rect 2828 37492 2884 37502
rect 2828 37398 2884 37436
rect 2716 36652 2884 36708
rect 2492 36430 2494 36482
rect 2546 36430 2548 36482
rect 2268 35758 2270 35810
rect 2322 35758 2324 35810
rect 2268 35746 2324 35758
rect 2380 36372 2436 36382
rect 2380 35364 2436 36316
rect 2492 35922 2548 36430
rect 2716 36484 2772 36494
rect 2716 36390 2772 36428
rect 2828 36148 2884 36652
rect 3052 36260 3108 37996
rect 3164 37380 3220 40572
rect 3276 37492 3332 40684
rect 3388 40402 3444 40414
rect 3388 40350 3390 40402
rect 3442 40350 3444 40402
rect 3388 40292 3444 40350
rect 3388 40226 3444 40236
rect 3612 40402 3668 43260
rect 3724 43250 3780 43260
rect 3612 40350 3614 40402
rect 3666 40350 3668 40402
rect 3612 40292 3668 40350
rect 3612 40226 3668 40236
rect 3948 39620 4004 45276
rect 4060 45266 4116 45276
rect 4172 45106 4228 45388
rect 4172 45054 4174 45106
rect 4226 45054 4228 45106
rect 4172 45042 4228 45054
rect 4476 44716 4740 44726
rect 4532 44660 4580 44716
rect 4636 44660 4684 44716
rect 4476 44650 4740 44660
rect 5740 44212 5796 44222
rect 5404 44210 5796 44212
rect 5404 44158 5742 44210
rect 5794 44158 5796 44210
rect 5404 44156 5796 44158
rect 4844 43652 4900 43662
rect 4844 43538 4900 43596
rect 5292 43652 5348 43662
rect 5292 43558 5348 43596
rect 4844 43486 4846 43538
rect 4898 43486 4900 43538
rect 4844 43474 4900 43486
rect 4060 43428 4116 43438
rect 4060 43334 4116 43372
rect 4508 43426 4564 43438
rect 4508 43374 4510 43426
rect 4562 43374 4564 43426
rect 4508 43316 4564 43374
rect 4508 43250 4564 43260
rect 4476 43148 4740 43158
rect 4532 43092 4580 43148
rect 4636 43092 4684 43148
rect 4476 43082 4740 43092
rect 5292 41972 5348 41982
rect 5404 41972 5460 44156
rect 5740 44146 5796 44156
rect 5852 43426 5908 43438
rect 5852 43374 5854 43426
rect 5906 43374 5908 43426
rect 5852 42308 5908 43374
rect 5852 42242 5908 42252
rect 5292 41970 5796 41972
rect 5292 41918 5294 41970
rect 5346 41918 5796 41970
rect 5292 41916 5796 41918
rect 5292 41906 5348 41916
rect 4060 41860 4116 41870
rect 4060 41766 4116 41804
rect 4476 41580 4740 41590
rect 4532 41524 4580 41580
rect 4636 41524 4684 41580
rect 4476 41514 4740 41524
rect 3948 39526 4004 39564
rect 4060 41188 4116 41198
rect 3388 39506 3444 39518
rect 3388 39454 3390 39506
rect 3442 39454 3444 39506
rect 3388 39284 3444 39454
rect 3500 39396 3556 39406
rect 3500 39302 3556 39340
rect 3388 38948 3444 39228
rect 3612 39060 3668 39070
rect 3500 38948 3556 38958
rect 3388 38892 3500 38948
rect 3500 38854 3556 38892
rect 3612 38050 3668 39004
rect 3836 38836 3892 38846
rect 3836 38742 3892 38780
rect 3612 37998 3614 38050
rect 3666 37998 3668 38050
rect 3612 37604 3668 37998
rect 3612 37538 3668 37548
rect 3836 38388 3892 38398
rect 3276 37436 3444 37492
rect 3164 37324 3332 37380
rect 3164 37156 3220 37166
rect 3164 37062 3220 37100
rect 3276 36932 3332 37324
rect 3164 36876 3332 36932
rect 3164 36596 3220 36876
rect 3164 36530 3220 36540
rect 3276 36484 3332 36494
rect 3276 36390 3332 36428
rect 3052 36204 3332 36260
rect 2828 36082 2884 36092
rect 2492 35870 2494 35922
rect 2546 35870 2548 35922
rect 2492 35858 2548 35870
rect 2716 35812 2772 35822
rect 2604 35700 2660 35710
rect 2604 35606 2660 35644
rect 2716 35698 2772 35756
rect 2940 35756 3220 35812
rect 2716 35646 2718 35698
rect 2770 35646 2772 35698
rect 2716 35634 2772 35646
rect 2828 35698 2884 35710
rect 2828 35646 2830 35698
rect 2882 35646 2884 35698
rect 2828 35364 2884 35646
rect 2380 35308 2884 35364
rect 2156 34850 2212 34860
rect 2268 34802 2324 34814
rect 2268 34750 2270 34802
rect 2322 34750 2324 34802
rect 2044 34412 2212 34468
rect 2044 34244 2100 34254
rect 2044 34150 2100 34188
rect 2044 33124 2100 33134
rect 2044 33030 2100 33068
rect 2044 31220 2100 31230
rect 1932 31164 2044 31220
rect 2044 31154 2100 31164
rect 2044 30996 2100 31006
rect 1932 30994 2100 30996
rect 1932 30942 2046 30994
rect 2098 30942 2100 30994
rect 1932 30940 2100 30942
rect 1708 30772 1764 30782
rect 1708 30212 1764 30716
rect 1708 30210 1876 30212
rect 1708 30158 1710 30210
rect 1762 30158 1876 30210
rect 1708 30156 1876 30158
rect 1708 30146 1764 30156
rect 1820 29650 1876 30156
rect 1820 29598 1822 29650
rect 1874 29598 1876 29650
rect 1820 29586 1876 29598
rect 1484 28242 1540 28252
rect 1820 28420 1876 28430
rect 1708 27858 1764 27870
rect 1708 27806 1710 27858
rect 1762 27806 1764 27858
rect 1708 27748 1764 27806
rect 1708 27188 1764 27692
rect 1708 27122 1764 27132
rect 1708 25396 1764 25406
rect 1708 25302 1764 25340
rect 1484 25060 1540 25070
rect 1484 8428 1540 25004
rect 1708 23826 1764 23838
rect 1708 23774 1710 23826
rect 1762 23774 1764 23826
rect 1708 23604 1764 23774
rect 1708 23538 1764 23548
rect 1708 22258 1764 22270
rect 1708 22206 1710 22258
rect 1762 22206 1764 22258
rect 1708 21812 1764 22206
rect 1708 21746 1764 21756
rect 1708 20578 1764 20590
rect 1708 20526 1710 20578
rect 1762 20526 1764 20578
rect 1708 20020 1764 20526
rect 1708 19954 1764 19964
rect 1708 18450 1764 18462
rect 1708 18398 1710 18450
rect 1762 18398 1764 18450
rect 1708 18228 1764 18398
rect 1708 18162 1764 18172
rect 1708 16882 1764 16894
rect 1708 16830 1710 16882
rect 1762 16830 1764 16882
rect 1708 16436 1764 16830
rect 1708 16370 1764 16380
rect 1820 15540 1876 28364
rect 1932 22260 1988 30940
rect 2044 30930 2100 30940
rect 2044 30100 2100 30110
rect 2044 30006 2100 30044
rect 2044 28532 2100 28542
rect 2044 28082 2100 28476
rect 2044 28030 2046 28082
rect 2098 28030 2100 28082
rect 2044 28018 2100 28030
rect 2044 25396 2100 25406
rect 2156 25396 2212 34412
rect 2268 33348 2324 34750
rect 2492 34692 2548 35308
rect 2828 35028 2884 35038
rect 2940 35028 2996 35756
rect 3164 35698 3220 35756
rect 3164 35646 3166 35698
rect 3218 35646 3220 35698
rect 3164 35634 3220 35646
rect 2828 35026 2996 35028
rect 2828 34974 2830 35026
rect 2882 34974 2996 35026
rect 2828 34972 2996 34974
rect 3052 35588 3108 35598
rect 2828 34962 2884 34972
rect 2604 34916 2660 34926
rect 2660 34860 2772 34916
rect 2604 34850 2660 34860
rect 2716 34802 2772 34860
rect 2716 34750 2718 34802
rect 2770 34750 2772 34802
rect 2716 34738 2772 34750
rect 2828 34804 2884 34814
rect 2828 34802 2996 34804
rect 2828 34750 2830 34802
rect 2882 34750 2996 34802
rect 2828 34748 2996 34750
rect 2828 34738 2884 34748
rect 2940 34692 2996 34748
rect 2492 34690 2660 34692
rect 2492 34638 2494 34690
rect 2546 34638 2660 34690
rect 2492 34636 2660 34638
rect 2492 34626 2548 34636
rect 2268 33282 2324 33292
rect 2492 34018 2548 34030
rect 2492 33966 2494 34018
rect 2546 33966 2548 34018
rect 2492 33236 2548 33966
rect 2492 33170 2548 33180
rect 2604 33346 2660 34636
rect 2940 34626 2996 34636
rect 2828 34580 2884 34590
rect 2604 33294 2606 33346
rect 2658 33294 2660 33346
rect 2604 32900 2660 33294
rect 2268 32844 2660 32900
rect 2716 34524 2828 34580
rect 2268 31218 2324 32844
rect 2268 31166 2270 31218
rect 2322 31166 2324 31218
rect 2268 31154 2324 31166
rect 2716 31108 2772 34524
rect 2828 34514 2884 34524
rect 3052 33572 3108 35532
rect 3276 35476 3332 36204
rect 3388 35924 3444 37436
rect 3612 37268 3668 37278
rect 3612 36594 3668 37212
rect 3612 36542 3614 36594
rect 3666 36542 3668 36594
rect 3612 36530 3668 36542
rect 3836 36372 3892 38332
rect 3948 38164 4004 38174
rect 3948 38070 4004 38108
rect 4060 37938 4116 41132
rect 5740 41188 5796 41916
rect 5852 41188 5908 41198
rect 5740 41186 5908 41188
rect 5740 41134 5854 41186
rect 5906 41134 5908 41186
rect 5740 41132 5908 41134
rect 4172 40516 4228 40526
rect 4956 40516 5012 40526
rect 4172 40514 4340 40516
rect 4172 40462 4174 40514
rect 4226 40462 4340 40514
rect 4172 40460 4340 40462
rect 4172 40450 4228 40460
rect 4284 38836 4340 40460
rect 4476 40012 4740 40022
rect 4532 39956 4580 40012
rect 4636 39956 4684 40012
rect 4476 39946 4740 39956
rect 4956 39506 5012 40460
rect 5068 40404 5124 40414
rect 5068 39618 5124 40348
rect 5740 40404 5796 41132
rect 5852 41122 5908 41132
rect 5740 40310 5796 40348
rect 5404 40292 5460 40302
rect 5068 39566 5070 39618
rect 5122 39566 5124 39618
rect 5068 39554 5124 39566
rect 5180 40290 5460 40292
rect 5180 40238 5406 40290
rect 5458 40238 5460 40290
rect 5180 40236 5460 40238
rect 4956 39454 4958 39506
rect 5010 39454 5012 39506
rect 4956 39442 5012 39454
rect 4284 38742 4340 38780
rect 4476 38444 4740 38454
rect 4532 38388 4580 38444
rect 4636 38388 4684 38444
rect 4476 38378 4740 38388
rect 4956 38276 5012 38286
rect 4956 38182 5012 38220
rect 4732 38052 4788 38062
rect 4732 37958 4788 37996
rect 4060 37886 4062 37938
rect 4114 37886 4116 37938
rect 4060 37874 4116 37886
rect 4284 37938 4340 37950
rect 4284 37886 4286 37938
rect 4338 37886 4340 37938
rect 3612 36370 3892 36372
rect 3612 36318 3838 36370
rect 3890 36318 3892 36370
rect 3612 36316 3892 36318
rect 3500 35924 3556 35934
rect 3388 35922 3556 35924
rect 3388 35870 3502 35922
rect 3554 35870 3556 35922
rect 3388 35868 3556 35870
rect 3500 35858 3556 35868
rect 3500 35588 3556 35598
rect 3500 35494 3556 35532
rect 3164 35420 3332 35476
rect 3164 34692 3220 35420
rect 3612 35308 3668 36316
rect 3836 36306 3892 36316
rect 3948 37604 4004 37614
rect 3948 36148 4004 37548
rect 4284 36484 4340 37886
rect 4476 36876 4740 36886
rect 4532 36820 4580 36876
rect 4636 36820 4684 36876
rect 4476 36810 4740 36820
rect 3836 36092 4004 36148
rect 4060 36428 4340 36484
rect 3164 34626 3220 34636
rect 3276 35252 3668 35308
rect 3724 35810 3780 35822
rect 3724 35758 3726 35810
rect 3778 35758 3780 35810
rect 3052 33506 3108 33516
rect 2604 31052 2772 31108
rect 2828 33348 2884 33358
rect 2380 30098 2436 30110
rect 2380 30046 2382 30098
rect 2434 30046 2436 30098
rect 2380 29988 2436 30046
rect 2044 25394 2212 25396
rect 2044 25342 2046 25394
rect 2098 25342 2212 25394
rect 2044 25340 2212 25342
rect 2268 29426 2324 29438
rect 2268 29374 2270 29426
rect 2322 29374 2324 29426
rect 2044 25330 2100 25340
rect 2268 25284 2324 29374
rect 2380 28980 2436 29932
rect 2380 28914 2436 28924
rect 2604 28754 2660 31052
rect 2604 28702 2606 28754
rect 2658 28702 2660 28754
rect 2604 28690 2660 28702
rect 2716 29986 2772 29998
rect 2716 29934 2718 29986
rect 2770 29934 2772 29986
rect 2380 28644 2436 28654
rect 2716 28644 2772 29934
rect 2828 29316 2884 33292
rect 3164 33236 3220 33246
rect 3164 33142 3220 33180
rect 3276 32788 3332 35252
rect 3388 34018 3444 34030
rect 3388 33966 3390 34018
rect 3442 33966 3444 34018
rect 3388 33236 3444 33966
rect 3500 33236 3556 33246
rect 3388 33234 3556 33236
rect 3388 33182 3502 33234
rect 3554 33182 3556 33234
rect 3388 33180 3556 33182
rect 3164 32732 3332 32788
rect 2940 32564 2996 32574
rect 2940 32562 3108 32564
rect 2940 32510 2942 32562
rect 2994 32510 3108 32562
rect 2940 32508 3108 32510
rect 2940 32498 2996 32508
rect 2828 29250 2884 29260
rect 2940 31892 2996 31902
rect 2828 28644 2884 28654
rect 2716 28642 2884 28644
rect 2716 28590 2830 28642
rect 2882 28590 2884 28642
rect 2716 28588 2884 28590
rect 2380 28550 2436 28588
rect 2828 28578 2884 28588
rect 2940 28644 2996 31836
rect 3052 31332 3108 32508
rect 3164 31780 3220 32732
rect 3276 32562 3332 32574
rect 3276 32510 3278 32562
rect 3330 32510 3332 32562
rect 3276 31948 3332 32510
rect 3276 31892 3444 31948
rect 3276 31780 3332 31790
rect 3164 31778 3332 31780
rect 3164 31726 3278 31778
rect 3330 31726 3332 31778
rect 3164 31724 3332 31726
rect 3276 31714 3332 31724
rect 3388 31780 3444 31892
rect 3052 31276 3220 31332
rect 3052 31108 3108 31118
rect 3052 31014 3108 31052
rect 3164 30212 3220 31276
rect 3388 31108 3444 31724
rect 3500 31444 3556 33180
rect 3612 33124 3668 33134
rect 3612 33030 3668 33068
rect 3612 32562 3668 32574
rect 3612 32510 3614 32562
rect 3666 32510 3668 32562
rect 3612 31892 3668 32510
rect 3724 32116 3780 35758
rect 3836 34354 3892 36092
rect 3836 34302 3838 34354
rect 3890 34302 3892 34354
rect 3836 34290 3892 34302
rect 3948 35476 4004 35486
rect 3836 33348 3892 33358
rect 3948 33348 4004 35420
rect 3836 33346 4004 33348
rect 3836 33294 3838 33346
rect 3890 33294 4004 33346
rect 3836 33292 4004 33294
rect 3836 33282 3892 33292
rect 4060 32340 4116 36428
rect 4284 36260 4340 36270
rect 4844 36260 4900 36270
rect 4284 36258 4900 36260
rect 4284 36206 4286 36258
rect 4338 36206 4846 36258
rect 4898 36206 4900 36258
rect 4284 36204 4900 36206
rect 4284 36194 4340 36204
rect 4284 36036 4340 36046
rect 4284 35588 4340 35980
rect 4620 35924 4676 35934
rect 4620 35830 4676 35868
rect 4284 35522 4340 35532
rect 4844 35364 4900 36204
rect 4476 35308 4740 35318
rect 4532 35252 4580 35308
rect 4636 35252 4684 35308
rect 4844 35298 4900 35308
rect 4476 35242 4740 35252
rect 4396 34356 4452 34366
rect 4284 34300 4396 34356
rect 4284 33572 4340 34300
rect 4396 34290 4452 34300
rect 4476 33740 4740 33750
rect 4532 33684 4580 33740
rect 4636 33684 4684 33740
rect 4476 33674 4740 33684
rect 4620 33572 4676 33582
rect 4284 33516 4452 33572
rect 4396 33346 4452 33516
rect 4396 33294 4398 33346
rect 4450 33294 4452 33346
rect 4396 33282 4452 33294
rect 4620 33346 4676 33516
rect 4620 33294 4622 33346
rect 4674 33294 4676 33346
rect 4620 33282 4676 33294
rect 5068 33348 5124 33358
rect 5068 33254 5124 33292
rect 3724 32050 3780 32060
rect 3948 32284 4116 32340
rect 4284 33236 4340 33246
rect 3612 31826 3668 31836
rect 3724 31890 3780 31902
rect 3724 31838 3726 31890
rect 3778 31838 3780 31890
rect 3724 31780 3780 31838
rect 3724 31714 3780 31724
rect 3500 31388 3668 31444
rect 2940 28578 2996 28588
rect 3052 30156 3220 30212
rect 3276 31052 3444 31108
rect 2492 28420 2548 28430
rect 2492 28326 2548 28364
rect 2716 28420 2772 28430
rect 2716 28326 2772 28364
rect 2492 27748 2548 27758
rect 2492 27654 2548 27692
rect 3052 26908 3108 30156
rect 3164 29988 3220 29998
rect 3164 29894 3220 29932
rect 3164 29540 3220 29550
rect 3276 29540 3332 31052
rect 3500 30996 3556 31006
rect 3612 30996 3668 31388
rect 3948 30996 4004 32284
rect 3500 30994 3668 30996
rect 3500 30942 3502 30994
rect 3554 30942 3668 30994
rect 3500 30940 3668 30942
rect 3500 30930 3556 30940
rect 3388 30884 3444 30894
rect 3388 30790 3444 30828
rect 3612 29876 3668 30940
rect 3836 30940 4004 30996
rect 4060 32116 4116 32126
rect 3724 29876 3780 29886
rect 3612 29820 3724 29876
rect 3724 29810 3780 29820
rect 3164 29538 3556 29540
rect 3164 29486 3166 29538
rect 3218 29486 3556 29538
rect 3164 29484 3556 29486
rect 3164 29474 3220 29484
rect 2940 26852 3108 26908
rect 3164 29316 3220 29326
rect 2940 26292 2996 26852
rect 2604 26236 2996 26292
rect 2492 25396 2548 25406
rect 2492 25302 2548 25340
rect 2156 25228 2324 25284
rect 2044 23828 2100 23838
rect 2044 23734 2100 23772
rect 2044 22260 2100 22270
rect 1932 22258 2100 22260
rect 1932 22206 2046 22258
rect 2098 22206 2100 22258
rect 1932 22204 2100 22206
rect 2044 22194 2100 22204
rect 2156 22036 2212 25228
rect 2604 23940 2660 26236
rect 1932 21980 2212 22036
rect 2268 23884 2660 23940
rect 1932 17108 1988 21980
rect 2268 21924 2324 23884
rect 3164 23828 3220 29260
rect 3276 28532 3332 28542
rect 3276 28438 3332 28476
rect 3500 28420 3556 29484
rect 3836 28754 3892 30940
rect 3836 28702 3838 28754
rect 3890 28702 3892 28754
rect 3836 28690 3892 28702
rect 3948 28644 4004 28654
rect 3948 28550 4004 28588
rect 3500 28326 3556 28364
rect 3724 28418 3780 28430
rect 3724 28366 3726 28418
rect 3778 28366 3780 28418
rect 3724 28196 3780 28366
rect 3724 28140 3892 28196
rect 3724 27972 3780 27982
rect 3500 27970 3780 27972
rect 3500 27918 3726 27970
rect 3778 27918 3780 27970
rect 3500 27916 3780 27918
rect 3388 27748 3444 27758
rect 3500 27748 3556 27916
rect 3724 27906 3780 27916
rect 3388 27746 3556 27748
rect 3388 27694 3390 27746
rect 3442 27694 3556 27746
rect 3388 27692 3556 27694
rect 3388 26964 3444 27692
rect 3388 26898 3444 26908
rect 3164 23762 3220 23772
rect 2492 23714 2548 23726
rect 2492 23662 2494 23714
rect 2546 23662 2548 23714
rect 2492 23604 2548 23662
rect 2492 23538 2548 23548
rect 2044 21868 2324 21924
rect 2380 23492 2436 23502
rect 2044 20690 2100 21868
rect 2380 21588 2436 23436
rect 2492 22146 2548 22158
rect 2492 22094 2494 22146
rect 2546 22094 2548 22146
rect 2492 21812 2548 22094
rect 2492 21746 2548 21756
rect 2380 21532 2548 21588
rect 2492 21364 2548 21532
rect 2044 20638 2046 20690
rect 2098 20638 2100 20690
rect 2044 20626 2100 20638
rect 2268 21308 2548 21364
rect 2268 20188 2324 21308
rect 2044 20132 2324 20188
rect 2492 20578 2548 20590
rect 2492 20526 2494 20578
rect 2546 20526 2548 20578
rect 2044 18674 2100 20132
rect 2492 20020 2548 20526
rect 2492 19954 2548 19964
rect 2044 18622 2046 18674
rect 2098 18622 2100 18674
rect 2044 18610 2100 18622
rect 2492 18338 2548 18350
rect 2492 18286 2494 18338
rect 2546 18286 2548 18338
rect 2492 18228 2548 18286
rect 2492 18162 2548 18172
rect 2044 17108 2100 17118
rect 1932 17106 2100 17108
rect 1932 17054 2046 17106
rect 2098 17054 2100 17106
rect 1932 17052 2100 17054
rect 2044 17042 2100 17052
rect 2492 16882 2548 16894
rect 2492 16830 2494 16882
rect 2546 16830 2548 16882
rect 2492 16436 2548 16830
rect 2492 16370 2548 16380
rect 2044 15540 2100 15550
rect 1820 15538 2100 15540
rect 1820 15486 2046 15538
rect 2098 15486 2100 15538
rect 1820 15484 2100 15486
rect 2044 15474 2100 15484
rect 1708 15314 1764 15326
rect 1708 15262 1710 15314
rect 1762 15262 1764 15314
rect 1708 14644 1764 15262
rect 1820 15204 1876 15214
rect 1876 15148 1988 15204
rect 1820 15138 1876 15148
rect 1708 14578 1764 14588
rect 1708 12852 1764 12862
rect 1708 12758 1764 12796
rect 1708 11282 1764 11294
rect 1708 11230 1710 11282
rect 1762 11230 1764 11282
rect 1708 11060 1764 11230
rect 1708 10994 1764 11004
rect 1708 9714 1764 9726
rect 1708 9662 1710 9714
rect 1762 9662 1764 9714
rect 1708 9268 1764 9662
rect 1932 9716 1988 15148
rect 2492 15202 2548 15214
rect 2492 15150 2494 15202
rect 2546 15150 2548 15202
rect 2492 14644 2548 15150
rect 2492 14578 2548 14588
rect 2044 13412 2100 13422
rect 2044 12850 2100 13356
rect 3836 13412 3892 28140
rect 3948 28084 4004 28094
rect 3948 27990 4004 28028
rect 3948 27748 4004 27758
rect 4060 27748 4116 32060
rect 4284 31778 4340 33180
rect 4508 33234 4564 33246
rect 4508 33182 4510 33234
rect 4562 33182 4564 33234
rect 4508 32340 4564 33182
rect 5180 33236 5236 40236
rect 5404 40226 5460 40236
rect 5628 40292 5684 40302
rect 5292 39620 5348 39630
rect 5292 39058 5348 39564
rect 5292 39006 5294 39058
rect 5346 39006 5348 39058
rect 5292 38994 5348 39006
rect 5628 38834 5684 40236
rect 5740 39508 5796 39518
rect 5740 38948 5796 39452
rect 5852 39060 5908 39070
rect 5852 38966 5908 39004
rect 5740 38854 5796 38892
rect 5628 38782 5630 38834
rect 5682 38782 5684 38834
rect 5628 38770 5684 38782
rect 5964 38668 6020 46510
rect 6076 40516 6132 48078
rect 6412 47572 6468 49534
rect 6524 49026 6580 49038
rect 6524 48974 6526 49026
rect 6578 48974 6580 49026
rect 6524 48356 6580 48974
rect 6636 49028 6692 49756
rect 7084 50034 7140 50046
rect 7084 49982 7086 50034
rect 7138 49982 7140 50034
rect 6972 49028 7028 49038
rect 6636 49026 7028 49028
rect 6636 48974 6974 49026
rect 7026 48974 7028 49026
rect 6636 48972 7028 48974
rect 6972 48962 7028 48972
rect 7084 48580 7140 49982
rect 7196 49924 7252 50764
rect 7308 50726 7364 50764
rect 7644 50370 7700 50382
rect 7644 50318 7646 50370
rect 7698 50318 7700 50370
rect 7532 49924 7588 49934
rect 7196 49922 7588 49924
rect 7196 49870 7198 49922
rect 7250 49870 7534 49922
rect 7586 49870 7588 49922
rect 7196 49868 7588 49870
rect 7196 49858 7252 49868
rect 7532 49858 7588 49868
rect 7420 48916 7476 48926
rect 6972 48524 7140 48580
rect 7308 48860 7420 48916
rect 6636 48356 6692 48366
rect 6524 48300 6636 48356
rect 6412 47506 6468 47516
rect 6636 48242 6692 48300
rect 6636 48190 6638 48242
rect 6690 48190 6692 48242
rect 6636 47458 6692 48190
rect 6636 47406 6638 47458
rect 6690 47406 6692 47458
rect 6188 47346 6244 47358
rect 6188 47294 6190 47346
rect 6242 47294 6244 47346
rect 6188 45556 6244 47294
rect 6412 46788 6468 46798
rect 6636 46788 6692 47406
rect 6412 46786 6692 46788
rect 6412 46734 6414 46786
rect 6466 46734 6692 46786
rect 6412 46732 6692 46734
rect 6412 46722 6468 46732
rect 6972 46676 7028 48524
rect 7084 48356 7140 48366
rect 7084 48262 7140 48300
rect 7196 48356 7252 48366
rect 7308 48356 7364 48860
rect 7420 48850 7476 48860
rect 7196 48354 7364 48356
rect 7196 48302 7198 48354
rect 7250 48302 7364 48354
rect 7196 48300 7364 48302
rect 7196 48290 7252 48300
rect 6748 46674 7028 46676
rect 6748 46622 6974 46674
rect 7026 46622 7028 46674
rect 6748 46620 7028 46622
rect 6188 45490 6244 45500
rect 6524 45778 6580 45790
rect 6524 45726 6526 45778
rect 6578 45726 6580 45778
rect 6524 45444 6580 45726
rect 6524 45378 6580 45388
rect 6636 45666 6692 45678
rect 6636 45614 6638 45666
rect 6690 45614 6692 45666
rect 6636 44548 6692 45614
rect 6748 45668 6804 46620
rect 6972 46610 7028 46620
rect 7084 48018 7140 48030
rect 7084 47966 7086 48018
rect 7138 47966 7140 48018
rect 6860 45892 6916 45902
rect 7084 45892 7140 47966
rect 7308 47458 7364 48300
rect 7308 47406 7310 47458
rect 7362 47406 7364 47458
rect 7308 47394 7364 47406
rect 7308 47124 7364 47134
rect 7308 46674 7364 47068
rect 7308 46622 7310 46674
rect 7362 46622 7364 46674
rect 7308 46610 7364 46622
rect 7532 46676 7588 46686
rect 6860 45890 7140 45892
rect 6860 45838 6862 45890
rect 6914 45838 7140 45890
rect 6860 45836 7140 45838
rect 6860 45826 6916 45836
rect 7084 45668 7140 45836
rect 6748 45612 6916 45668
rect 6748 45444 6804 45454
rect 6748 44994 6804 45388
rect 6748 44942 6750 44994
rect 6802 44942 6804 44994
rect 6748 44930 6804 44942
rect 6860 45106 6916 45612
rect 7084 45602 7140 45612
rect 7308 46002 7364 46014
rect 7308 45950 7310 46002
rect 7362 45950 7364 46002
rect 6860 45054 6862 45106
rect 6914 45054 6916 45106
rect 6300 44492 6692 44548
rect 6188 40516 6244 40526
rect 6076 40460 6188 40516
rect 6188 40422 6244 40460
rect 6076 39394 6132 39406
rect 6076 39342 6078 39394
rect 6130 39342 6132 39394
rect 6076 38948 6132 39342
rect 6076 38882 6132 38892
rect 6300 38668 6356 44492
rect 6860 44322 6916 45054
rect 6972 45556 7028 45566
rect 6972 45108 7028 45500
rect 6972 45106 7252 45108
rect 6972 45054 6974 45106
rect 7026 45054 7252 45106
rect 6972 45052 7252 45054
rect 6972 45042 7028 45052
rect 6860 44270 6862 44322
rect 6914 44270 6916 44322
rect 6860 44212 6916 44270
rect 6860 44146 6916 44156
rect 6860 43764 6916 43774
rect 6524 43652 6580 43662
rect 6524 43558 6580 43596
rect 6860 43538 6916 43708
rect 6860 43486 6862 43538
rect 6914 43486 6916 43538
rect 6860 43474 6916 43486
rect 7196 43762 7252 45052
rect 7196 43710 7198 43762
rect 7250 43710 7252 43762
rect 6860 43314 6916 43326
rect 6860 43262 6862 43314
rect 6914 43262 6916 43314
rect 6636 42308 6692 42318
rect 6524 42252 6636 42308
rect 6412 42084 6468 42094
rect 6412 41990 6468 42028
rect 6412 41076 6468 41086
rect 6524 41076 6580 42252
rect 6636 42242 6692 42252
rect 6412 41074 6580 41076
rect 6412 41022 6414 41074
rect 6466 41022 6580 41074
rect 6412 41020 6580 41022
rect 6412 41010 6468 41020
rect 5740 38612 6020 38668
rect 6188 38612 6356 38668
rect 6412 39620 6468 39630
rect 6412 38724 6468 39564
rect 5628 38050 5684 38062
rect 5628 37998 5630 38050
rect 5682 37998 5684 38050
rect 5628 37828 5684 37998
rect 5628 37762 5684 37772
rect 5740 36482 5796 38612
rect 5740 36430 5742 36482
rect 5794 36430 5796 36482
rect 5628 36372 5684 36382
rect 5516 36316 5628 36372
rect 5404 35588 5460 35598
rect 5180 33170 5236 33180
rect 5292 34692 5348 34702
rect 5292 32676 5348 34636
rect 5404 34356 5460 35532
rect 5404 34262 5460 34300
rect 5404 32676 5460 32686
rect 5292 32674 5460 32676
rect 5292 32622 5406 32674
rect 5458 32622 5460 32674
rect 5292 32620 5460 32622
rect 5404 32610 5460 32620
rect 4956 32564 5012 32574
rect 4956 32470 5012 32508
rect 4508 32284 4900 32340
rect 4476 32172 4740 32182
rect 4532 32116 4580 32172
rect 4636 32116 4684 32172
rect 4476 32106 4740 32116
rect 4284 31726 4286 31778
rect 4338 31726 4340 31778
rect 4284 31714 4340 31726
rect 4396 31106 4452 31118
rect 4396 31054 4398 31106
rect 4450 31054 4452 31106
rect 4396 30884 4452 31054
rect 4844 30996 4900 32284
rect 5516 31220 5572 36316
rect 5628 36306 5684 36316
rect 5740 35922 5796 36430
rect 6188 37826 6244 38612
rect 6412 38052 6468 38668
rect 6524 38668 6580 41020
rect 6748 41860 6804 41870
rect 6748 40404 6804 41804
rect 6748 39618 6804 40348
rect 6748 39566 6750 39618
rect 6802 39566 6804 39618
rect 6748 39554 6804 39566
rect 6748 38836 6804 38874
rect 6748 38770 6804 38780
rect 6860 38668 6916 43262
rect 7196 42084 7252 43710
rect 7308 43764 7364 45950
rect 7308 43698 7364 43708
rect 7532 42532 7588 46620
rect 7644 45892 7700 50318
rect 8092 49698 8148 49710
rect 8092 49646 8094 49698
rect 8146 49646 8148 49698
rect 8092 48916 8148 49646
rect 8204 49028 8260 55412
rect 10444 53506 10500 55412
rect 11788 55188 11844 55198
rect 11788 55094 11844 55132
rect 11900 55076 11956 55086
rect 12684 55076 12740 55412
rect 13692 55412 14420 55468
rect 16380 55412 16436 55422
rect 13580 55300 13636 55310
rect 13580 55206 13636 55244
rect 11900 55074 12516 55076
rect 11900 55022 11902 55074
rect 11954 55022 12516 55074
rect 11900 55020 12516 55022
rect 11900 55010 11956 55020
rect 12460 54852 12516 55020
rect 12684 55010 12740 55020
rect 12460 54796 13300 54852
rect 12460 54738 12516 54796
rect 12460 54686 12462 54738
rect 12514 54686 12516 54738
rect 12460 54674 12516 54686
rect 12796 54626 12852 54638
rect 12796 54574 12798 54626
rect 12850 54574 12852 54626
rect 12796 53844 12852 54574
rect 13244 54626 13300 54796
rect 13244 54574 13246 54626
rect 13298 54574 13300 54626
rect 13244 54562 13300 54574
rect 13692 54514 13748 55412
rect 16268 55410 16436 55412
rect 16268 55358 16382 55410
rect 16434 55358 16436 55410
rect 16268 55356 16436 55358
rect 14252 55188 14308 55198
rect 14252 55186 14868 55188
rect 14252 55134 14254 55186
rect 14306 55134 14868 55186
rect 14252 55132 14868 55134
rect 14252 55122 14308 55132
rect 14812 54738 14868 55132
rect 15820 54740 15876 54750
rect 14812 54686 14814 54738
rect 14866 54686 14868 54738
rect 14812 54674 14868 54686
rect 15260 54738 15876 54740
rect 15260 54686 15822 54738
rect 15874 54686 15876 54738
rect 15260 54684 15876 54686
rect 15260 54626 15316 54684
rect 15820 54674 15876 54684
rect 15260 54574 15262 54626
rect 15314 54574 15316 54626
rect 15260 54562 15316 54574
rect 13692 54462 13694 54514
rect 13746 54462 13748 54514
rect 13692 54450 13748 54462
rect 14588 54514 14644 54526
rect 14588 54462 14590 54514
rect 14642 54462 14644 54514
rect 12796 53778 12852 53788
rect 13804 54402 13860 54414
rect 13804 54350 13806 54402
rect 13858 54350 13860 54402
rect 10444 53454 10446 53506
rect 10498 53454 10500 53506
rect 9884 53060 9940 53070
rect 8764 52946 8820 52958
rect 8764 52894 8766 52946
rect 8818 52894 8820 52946
rect 8764 52164 8820 52894
rect 8988 52164 9044 52174
rect 8764 52162 9044 52164
rect 8764 52110 8990 52162
rect 9042 52110 9044 52162
rect 8764 52108 9044 52110
rect 9884 52164 9940 53004
rect 10220 52948 10276 52958
rect 10444 52948 10500 53454
rect 11564 53508 11620 53518
rect 10220 52946 10500 52948
rect 10220 52894 10222 52946
rect 10274 52894 10500 52946
rect 10220 52892 10500 52894
rect 10556 53060 10612 53070
rect 10220 52612 10276 52892
rect 10220 52546 10276 52556
rect 10444 52724 10500 52734
rect 10332 52500 10388 52510
rect 9996 52164 10052 52174
rect 9884 52162 10052 52164
rect 9884 52110 9998 52162
rect 10050 52110 10052 52162
rect 9884 52108 10052 52110
rect 8988 51940 9044 52108
rect 9996 52098 10052 52108
rect 10332 52162 10388 52444
rect 10444 52386 10500 52668
rect 10444 52334 10446 52386
rect 10498 52334 10500 52386
rect 10444 52322 10500 52334
rect 10332 52110 10334 52162
rect 10386 52110 10388 52162
rect 10332 52098 10388 52110
rect 8988 51380 9044 51884
rect 10108 51938 10164 51950
rect 10108 51886 10110 51938
rect 10162 51886 10164 51938
rect 10108 51828 10164 51886
rect 10108 51762 10164 51772
rect 10556 51492 10612 53004
rect 11116 53060 11172 53070
rect 10668 52948 10724 52958
rect 10668 52854 10724 52892
rect 10892 52948 10948 52958
rect 10892 52854 10948 52892
rect 11004 52724 11060 52734
rect 10780 52162 10836 52174
rect 10780 52110 10782 52162
rect 10834 52110 10836 52162
rect 10668 51492 10724 51502
rect 10556 51490 10724 51492
rect 10556 51438 10670 51490
rect 10722 51438 10724 51490
rect 10556 51436 10724 51438
rect 10668 51426 10724 51436
rect 10780 51492 10836 52110
rect 10780 51426 10836 51436
rect 10892 51604 10948 51614
rect 10892 51490 10948 51548
rect 10892 51438 10894 51490
rect 10946 51438 10948 51490
rect 10892 51426 10948 51438
rect 11004 51380 11060 52668
rect 11116 52162 11172 53004
rect 11340 52948 11396 52958
rect 11564 52948 11620 53452
rect 12348 53172 12404 53182
rect 12012 53060 12068 53070
rect 11340 52946 11508 52948
rect 11340 52894 11342 52946
rect 11394 52894 11508 52946
rect 11340 52892 11508 52894
rect 11340 52882 11396 52892
rect 11116 52110 11118 52162
rect 11170 52110 11172 52162
rect 11116 52098 11172 52110
rect 11340 52164 11396 52174
rect 11340 52070 11396 52108
rect 11116 51380 11172 51390
rect 11004 51378 11172 51380
rect 11004 51326 11118 51378
rect 11170 51326 11172 51378
rect 11004 51324 11172 51326
rect 8988 51314 9044 51324
rect 11116 51314 11172 51324
rect 11228 51378 11284 51390
rect 11228 51326 11230 51378
rect 11282 51326 11284 51378
rect 10780 51266 10836 51278
rect 10780 51214 10782 51266
rect 10834 51214 10836 51266
rect 10780 49924 10836 51214
rect 11228 50428 11284 51326
rect 11452 50484 11508 52892
rect 11564 52882 11620 52892
rect 11676 53058 12068 53060
rect 11676 53006 12014 53058
rect 12066 53006 12068 53058
rect 11676 53004 12068 53006
rect 11676 52724 11732 53004
rect 12012 52994 12068 53004
rect 12348 53058 12404 53116
rect 12796 53172 12852 53182
rect 12796 53078 12852 53116
rect 13804 53172 13860 54350
rect 13804 53106 13860 53116
rect 12348 53006 12350 53058
rect 12402 53006 12404 53058
rect 12348 52994 12404 53006
rect 11676 52386 11732 52668
rect 12684 52612 12740 52622
rect 12012 52388 12068 52398
rect 11676 52334 11678 52386
rect 11730 52334 11732 52386
rect 11676 52322 11732 52334
rect 11900 52386 12068 52388
rect 11900 52334 12014 52386
rect 12066 52334 12068 52386
rect 11900 52332 12068 52334
rect 11900 52162 11956 52332
rect 12012 52322 12068 52332
rect 11900 52110 11902 52162
rect 11954 52110 11956 52162
rect 11900 52098 11956 52110
rect 12348 52164 12404 52174
rect 12348 52070 12404 52108
rect 11900 51938 11956 51950
rect 11900 51886 11902 51938
rect 11954 51886 11956 51938
rect 11116 50372 11284 50428
rect 11340 50428 11508 50484
rect 11564 51492 11620 51502
rect 11116 50036 11172 50372
rect 11340 50260 11396 50428
rect 11116 49970 11172 49980
rect 11228 50204 11396 50260
rect 10780 49858 10836 49868
rect 8204 48962 8260 48972
rect 8428 49810 8484 49822
rect 8428 49758 8430 49810
rect 8482 49758 8484 49810
rect 8092 48850 8148 48860
rect 8428 48916 8484 49758
rect 8988 49812 9044 49822
rect 8988 49718 9044 49756
rect 10556 49812 10612 49822
rect 11228 49812 11284 50204
rect 11564 50148 11620 51436
rect 11900 51268 11956 51886
rect 12012 51604 12068 51614
rect 12012 51510 12068 51548
rect 11900 51202 11956 51212
rect 12684 50428 12740 52556
rect 12796 52500 12852 52510
rect 12796 52274 12852 52444
rect 12796 52222 12798 52274
rect 12850 52222 12852 52274
rect 12796 52210 12852 52222
rect 13020 52386 13076 52398
rect 13020 52334 13022 52386
rect 13074 52334 13076 52386
rect 11900 50372 11956 50382
rect 11340 50092 11620 50148
rect 11676 50370 12180 50372
rect 11676 50318 11902 50370
rect 11954 50318 12180 50370
rect 11676 50316 12180 50318
rect 11340 50034 11396 50092
rect 11340 49982 11342 50034
rect 11394 49982 11396 50034
rect 11340 49970 11396 49982
rect 11564 49812 11620 49822
rect 11676 49812 11732 50316
rect 11900 50306 11956 50316
rect 12012 50036 12068 50046
rect 12124 50036 12180 50316
rect 12572 50370 12628 50382
rect 12684 50372 12964 50428
rect 12572 50318 12574 50370
rect 12626 50318 12628 50370
rect 12572 50036 12628 50318
rect 12124 49980 12572 50036
rect 12012 49942 12068 49980
rect 10612 49756 10724 49812
rect 11228 49756 11396 49812
rect 10556 49718 10612 49756
rect 8428 48850 8484 48860
rect 10108 49698 10164 49710
rect 10108 49646 10110 49698
rect 10162 49646 10164 49698
rect 10108 49252 10164 49646
rect 10556 49588 10612 49598
rect 9660 48802 9716 48814
rect 9660 48750 9662 48802
rect 9714 48750 9716 48802
rect 8316 48468 8372 48478
rect 7756 47570 7812 47582
rect 7756 47518 7758 47570
rect 7810 47518 7812 47570
rect 7756 46676 7812 47518
rect 8316 47458 8372 48412
rect 9660 48468 9716 48750
rect 9660 48402 9716 48412
rect 9660 48242 9716 48254
rect 9660 48190 9662 48242
rect 9714 48190 9716 48242
rect 8316 47406 8318 47458
rect 8370 47406 8372 47458
rect 8316 47124 8372 47406
rect 8764 47460 8820 47470
rect 8764 47366 8820 47404
rect 8316 47058 8372 47068
rect 9212 47348 9268 47358
rect 9660 47348 9716 48190
rect 9212 47346 9716 47348
rect 9212 47294 9214 47346
rect 9266 47294 9716 47346
rect 9212 47292 9716 47294
rect 8988 46900 9044 46910
rect 7868 46788 7924 46798
rect 7868 46694 7924 46732
rect 7756 46610 7812 46620
rect 8652 45892 8708 45902
rect 7644 45890 8260 45892
rect 7644 45838 7646 45890
rect 7698 45838 8260 45890
rect 7644 45836 8260 45838
rect 7644 45826 7700 45836
rect 8092 45668 8148 45678
rect 8092 45574 8148 45612
rect 7980 45444 8036 45454
rect 7980 45218 8036 45388
rect 8204 45330 8260 45836
rect 8652 45798 8708 45836
rect 8764 45780 8820 45790
rect 8820 45724 8932 45780
rect 8764 45714 8820 45724
rect 8204 45278 8206 45330
rect 8258 45278 8260 45330
rect 8204 45266 8260 45278
rect 8316 45668 8372 45678
rect 7980 45166 7982 45218
rect 8034 45166 8036 45218
rect 7980 45154 8036 45166
rect 7756 45108 7812 45118
rect 7756 45014 7812 45052
rect 8204 44994 8260 45006
rect 8204 44942 8206 44994
rect 8258 44942 8260 44994
rect 7980 44324 8036 44334
rect 7980 43764 8036 44268
rect 8092 44212 8148 44222
rect 8092 44118 8148 44156
rect 8204 43876 8260 44942
rect 7756 43652 7812 43662
rect 7756 43558 7812 43596
rect 7868 43428 7924 43438
rect 7868 42756 7924 43372
rect 7980 42866 8036 43708
rect 7980 42814 7982 42866
rect 8034 42814 8036 42866
rect 7980 42802 8036 42814
rect 8092 43820 8260 43876
rect 7196 42018 7252 42028
rect 7308 42476 7588 42532
rect 7756 42700 7868 42756
rect 7196 40516 7252 40526
rect 7196 39506 7252 40460
rect 7308 39620 7364 42476
rect 7756 42420 7812 42700
rect 7868 42662 7924 42700
rect 7420 42364 7812 42420
rect 7420 41970 7476 42364
rect 7420 41918 7422 41970
rect 7474 41918 7476 41970
rect 7420 41906 7476 41918
rect 7644 42084 7700 42094
rect 7644 41298 7700 42028
rect 7644 41246 7646 41298
rect 7698 41246 7700 41298
rect 7644 41234 7700 41246
rect 7868 40964 7924 40974
rect 7868 40962 8036 40964
rect 7868 40910 7870 40962
rect 7922 40910 8036 40962
rect 7868 40908 8036 40910
rect 7868 40898 7924 40908
rect 7756 39844 7812 39854
rect 7980 39844 8036 40908
rect 8092 40628 8148 43820
rect 8316 43204 8372 45612
rect 8540 44434 8596 44446
rect 8540 44382 8542 44434
rect 8594 44382 8596 44434
rect 8540 43764 8596 44382
rect 8316 43148 8484 43204
rect 8316 42978 8372 42990
rect 8316 42926 8318 42978
rect 8370 42926 8372 42978
rect 8316 42868 8372 42926
rect 8316 42802 8372 42812
rect 8204 42754 8260 42766
rect 8204 42702 8206 42754
rect 8258 42702 8260 42754
rect 8204 42644 8260 42702
rect 8428 42644 8484 43148
rect 8204 42578 8260 42588
rect 8316 42588 8484 42644
rect 8092 40572 8260 40628
rect 8092 40404 8148 40442
rect 8092 40338 8148 40348
rect 8204 40292 8260 40572
rect 8204 40226 8260 40236
rect 7364 39564 7588 39620
rect 7308 39554 7364 39564
rect 7196 39454 7198 39506
rect 7250 39454 7252 39506
rect 7196 39442 7252 39454
rect 7420 39060 7476 39070
rect 7308 38948 7364 38958
rect 7420 38948 7476 39004
rect 7308 38946 7476 38948
rect 7308 38894 7310 38946
rect 7362 38894 7476 38946
rect 7308 38892 7476 38894
rect 7308 38882 7364 38892
rect 6524 38612 6804 38668
rect 6860 38612 7028 38668
rect 6524 38052 6580 38062
rect 6412 38050 6580 38052
rect 6412 37998 6526 38050
rect 6578 37998 6580 38050
rect 6412 37996 6580 37998
rect 6188 37774 6190 37826
rect 6242 37774 6244 37826
rect 5964 36372 6020 36382
rect 5964 36278 6020 36316
rect 5740 35870 5742 35922
rect 5794 35870 5796 35922
rect 5740 35858 5796 35870
rect 5740 35364 5796 35374
rect 5628 34802 5684 34814
rect 5628 34750 5630 34802
rect 5682 34750 5684 34802
rect 5628 32004 5684 34750
rect 5628 31938 5684 31948
rect 5516 31154 5572 31164
rect 5628 31106 5684 31118
rect 5628 31054 5630 31106
rect 5682 31054 5684 31106
rect 5516 30996 5572 31006
rect 4844 30994 5012 30996
rect 4844 30942 4846 30994
rect 4898 30942 5012 30994
rect 4844 30940 5012 30942
rect 4844 30930 4900 30940
rect 4396 30818 4452 30828
rect 4476 30604 4740 30614
rect 4532 30548 4580 30604
rect 4636 30548 4684 30604
rect 4476 30538 4740 30548
rect 4956 30434 5012 30940
rect 5516 30902 5572 30940
rect 4956 30382 4958 30434
rect 5010 30382 5012 30434
rect 4956 30370 5012 30382
rect 5068 30098 5124 30110
rect 5068 30046 5070 30098
rect 5122 30046 5124 30098
rect 4172 29988 4228 29998
rect 4172 29894 4228 29932
rect 4620 29988 4676 29998
rect 4956 29988 5012 29998
rect 4620 29986 5012 29988
rect 4620 29934 4622 29986
rect 4674 29934 4958 29986
rect 5010 29934 5012 29986
rect 4620 29932 5012 29934
rect 4620 29922 4676 29932
rect 4620 29428 4676 29438
rect 4620 29334 4676 29372
rect 4476 29036 4740 29046
rect 4532 28980 4580 29036
rect 4636 28980 4684 29036
rect 4476 28970 4740 28980
rect 4396 28420 4452 28430
rect 3948 27746 4116 27748
rect 3948 27694 3950 27746
rect 4002 27694 4116 27746
rect 3948 27692 4116 27694
rect 4284 28418 4452 28420
rect 4284 28366 4398 28418
rect 4450 28366 4452 28418
rect 4284 28364 4452 28366
rect 4284 27858 4340 28364
rect 4396 28354 4452 28364
rect 4844 28308 4900 28318
rect 4844 28082 4900 28252
rect 4844 28030 4846 28082
rect 4898 28030 4900 28082
rect 4844 28018 4900 28030
rect 4956 27972 5012 29932
rect 5068 29988 5124 30046
rect 5068 29316 5124 29932
rect 5628 29540 5684 31054
rect 5740 29764 5796 35308
rect 6188 34916 6244 37774
rect 6300 37492 6356 37502
rect 6524 37492 6580 37996
rect 6748 37938 6804 38612
rect 6748 37886 6750 37938
rect 6802 37886 6804 37938
rect 6748 37874 6804 37886
rect 6300 37490 6580 37492
rect 6300 37438 6302 37490
rect 6354 37438 6580 37490
rect 6300 37436 6580 37438
rect 6860 37826 6916 37838
rect 6860 37774 6862 37826
rect 6914 37774 6916 37826
rect 6300 37426 6356 37436
rect 6748 36372 6804 36382
rect 6748 36278 6804 36316
rect 6300 35586 6356 35598
rect 6300 35534 6302 35586
rect 6354 35534 6356 35586
rect 6300 35140 6356 35534
rect 6300 35074 6356 35084
rect 6524 34916 6580 34926
rect 6188 34914 6580 34916
rect 6188 34862 6526 34914
rect 6578 34862 6580 34914
rect 6188 34860 6580 34862
rect 6524 34850 6580 34860
rect 6188 34692 6244 34702
rect 6188 34598 6244 34636
rect 6636 34356 6692 34366
rect 6636 34262 6692 34300
rect 6524 34244 6580 34254
rect 5852 34018 5908 34030
rect 5852 33966 5854 34018
rect 5906 33966 5908 34018
rect 5852 30996 5908 33966
rect 5964 33348 6020 33358
rect 5964 33254 6020 33292
rect 6524 32562 6580 34188
rect 6636 33572 6692 33582
rect 6636 32788 6692 33516
rect 6748 32788 6804 32798
rect 6636 32786 6804 32788
rect 6636 32734 6750 32786
rect 6802 32734 6804 32786
rect 6636 32732 6804 32734
rect 6748 32722 6804 32732
rect 6524 32510 6526 32562
rect 6578 32510 6580 32562
rect 6524 32498 6580 32510
rect 6636 32340 6692 32350
rect 6076 31332 6132 31342
rect 5964 30996 6020 31006
rect 5852 30940 5964 30996
rect 5964 30930 6020 30940
rect 5852 29988 5908 29998
rect 5852 29894 5908 29932
rect 5740 29708 5908 29764
rect 5852 29540 5908 29708
rect 6076 29652 6132 31276
rect 6300 30882 6356 30894
rect 6300 30830 6302 30882
rect 6354 30830 6356 30882
rect 6188 30100 6244 30110
rect 6188 30006 6244 30044
rect 6188 29652 6244 29662
rect 6076 29650 6244 29652
rect 6076 29598 6190 29650
rect 6242 29598 6244 29650
rect 6076 29596 6244 29598
rect 6188 29586 6244 29596
rect 5852 29484 6132 29540
rect 5628 29474 5684 29484
rect 5068 29250 5124 29260
rect 5740 29426 5796 29438
rect 5740 29374 5742 29426
rect 5794 29374 5796 29426
rect 5740 28644 5796 29374
rect 5740 28578 5796 28588
rect 5292 28532 5348 28542
rect 5292 28084 5348 28476
rect 5964 28420 6020 28430
rect 4956 27906 5012 27916
rect 5068 27970 5124 27982
rect 5068 27918 5070 27970
rect 5122 27918 5124 27970
rect 4284 27806 4286 27858
rect 4338 27806 4340 27858
rect 3948 27682 4004 27692
rect 4284 27636 4340 27806
rect 4284 27570 4340 27580
rect 4476 27468 4740 27478
rect 4532 27412 4580 27468
rect 4636 27412 4684 27468
rect 4476 27402 4740 27412
rect 4732 26962 4788 26974
rect 4732 26910 4734 26962
rect 4786 26910 4788 26962
rect 4732 26908 4788 26910
rect 5068 26908 5124 27918
rect 4732 26852 5124 26908
rect 4476 25900 4740 25910
rect 4532 25844 4580 25900
rect 4636 25844 4684 25900
rect 4476 25834 4740 25844
rect 4732 25060 4788 25070
rect 4844 25060 4900 26852
rect 5292 26292 5348 28028
rect 5852 28308 5908 28318
rect 5404 27860 5460 27870
rect 5404 27746 5460 27804
rect 5404 27694 5406 27746
rect 5458 27694 5460 27746
rect 5404 27682 5460 27694
rect 5516 27858 5572 27870
rect 5516 27806 5518 27858
rect 5570 27806 5572 27858
rect 5516 27748 5572 27806
rect 5852 27858 5908 28252
rect 5852 27806 5854 27858
rect 5906 27806 5908 27858
rect 5852 27794 5908 27806
rect 5516 27682 5572 27692
rect 5964 27748 6020 28364
rect 6076 28196 6132 29484
rect 6188 28642 6244 28654
rect 6188 28590 6190 28642
rect 6242 28590 6244 28642
rect 6188 28308 6244 28590
rect 6300 28644 6356 30830
rect 6636 30322 6692 32284
rect 6636 30270 6638 30322
rect 6690 30270 6692 30322
rect 6636 30258 6692 30270
rect 6860 30210 6916 37774
rect 6860 30158 6862 30210
rect 6914 30158 6916 30210
rect 6636 30100 6692 30110
rect 6636 30006 6692 30044
rect 6412 29986 6468 29998
rect 6412 29934 6414 29986
rect 6466 29934 6468 29986
rect 6412 29876 6468 29934
rect 6412 29810 6468 29820
rect 6412 29538 6468 29550
rect 6412 29486 6414 29538
rect 6466 29486 6468 29538
rect 6412 29428 6468 29486
rect 6412 29372 6692 29428
rect 6524 28644 6580 28654
rect 6300 28642 6580 28644
rect 6300 28590 6526 28642
rect 6578 28590 6580 28642
rect 6300 28588 6580 28590
rect 6524 28578 6580 28588
rect 6636 28308 6692 29372
rect 6188 28252 6692 28308
rect 6076 28140 6244 28196
rect 5964 27682 6020 27692
rect 6076 27970 6132 27982
rect 6076 27918 6078 27970
rect 6130 27918 6132 27970
rect 5964 27076 6020 27086
rect 5740 26964 5796 26974
rect 5516 26292 5572 26302
rect 5292 26290 5572 26292
rect 5292 26238 5518 26290
rect 5570 26238 5572 26290
rect 5292 26236 5572 26238
rect 5516 26226 5572 26236
rect 4788 25004 4900 25060
rect 4732 24994 4788 25004
rect 4476 24332 4740 24342
rect 4532 24276 4580 24332
rect 4636 24276 4684 24332
rect 4476 24266 4740 24276
rect 5740 23268 5796 26908
rect 5964 26292 6020 27020
rect 6076 26516 6132 27918
rect 6188 26908 6244 28140
rect 6412 27972 6468 27982
rect 6412 27186 6468 27916
rect 6412 27134 6414 27186
rect 6466 27134 6468 27186
rect 6412 27122 6468 27134
rect 6188 26852 6356 26908
rect 6076 26450 6132 26460
rect 5964 26198 6020 26236
rect 5852 23268 5908 23278
rect 5740 23212 5852 23268
rect 5852 23202 5908 23212
rect 4476 22764 4740 22774
rect 4532 22708 4580 22764
rect 4636 22708 4684 22764
rect 4476 22698 4740 22708
rect 4476 21196 4740 21206
rect 4532 21140 4580 21196
rect 4636 21140 4684 21196
rect 4476 21130 4740 21140
rect 4476 19628 4740 19638
rect 4532 19572 4580 19628
rect 4636 19572 4684 19628
rect 4476 19562 4740 19572
rect 4476 18060 4740 18070
rect 4532 18004 4580 18060
rect 4636 18004 4684 18060
rect 4476 17994 4740 18004
rect 4476 16492 4740 16502
rect 4532 16436 4580 16492
rect 4636 16436 4684 16492
rect 4476 16426 4740 16436
rect 4476 14924 4740 14934
rect 4532 14868 4580 14924
rect 4636 14868 4684 14924
rect 4476 14858 4740 14868
rect 3836 13346 3892 13356
rect 4476 13356 4740 13366
rect 4532 13300 4580 13356
rect 4636 13300 4684 13356
rect 4476 13290 4740 13300
rect 2044 12798 2046 12850
rect 2098 12798 2100 12850
rect 2044 12786 2100 12798
rect 2492 12852 2548 12862
rect 2492 12758 2548 12796
rect 4476 11788 4740 11798
rect 4532 11732 4580 11788
rect 4636 11732 4684 11788
rect 4476 11722 4740 11732
rect 2044 11284 2100 11294
rect 2044 11190 2100 11228
rect 6300 11284 6356 26852
rect 6300 11218 6356 11228
rect 2492 11170 2548 11182
rect 2492 11118 2494 11170
rect 2546 11118 2548 11170
rect 2492 11060 2548 11118
rect 2492 10994 2548 11004
rect 4476 10220 4740 10230
rect 4532 10164 4580 10220
rect 4636 10164 4684 10220
rect 4476 10154 4740 10164
rect 2380 10052 2436 10062
rect 2044 9716 2100 9726
rect 1932 9714 2100 9716
rect 1932 9662 2046 9714
rect 2098 9662 2100 9714
rect 1932 9660 2100 9662
rect 2044 9650 2100 9660
rect 1708 9202 1764 9212
rect 1484 8372 2100 8428
rect 1708 8146 1764 8158
rect 1708 8094 1710 8146
rect 1762 8094 1764 8146
rect 1708 8036 1764 8094
rect 2044 8146 2100 8372
rect 2044 8094 2046 8146
rect 2098 8094 2100 8146
rect 2044 8082 2100 8094
rect 1708 7476 1764 7980
rect 1708 7410 1764 7420
rect 1260 5842 1316 5852
rect 1708 5906 1764 5918
rect 1708 5854 1710 5906
rect 1762 5854 1764 5906
rect 1708 5684 1764 5854
rect 2156 5908 2212 5918
rect 2156 5794 2212 5852
rect 2156 5742 2158 5794
rect 2210 5742 2212 5794
rect 2156 5730 2212 5742
rect 1708 5236 1764 5628
rect 1820 5236 1876 5246
rect 1708 5234 1876 5236
rect 1708 5182 1822 5234
rect 1874 5182 1876 5234
rect 1708 5180 1876 5182
rect 1820 5170 1876 5180
rect 2044 4564 2100 4574
rect 2044 4470 2100 4508
rect 1708 4338 1764 4350
rect 1708 4286 1710 4338
rect 1762 4286 1764 4338
rect 1708 3892 1764 4286
rect 1708 3826 1764 3836
rect 2268 3668 2324 3678
rect 2380 3668 2436 9996
rect 6524 10052 6580 28252
rect 6748 27858 6804 27870
rect 6748 27806 6750 27858
rect 6802 27806 6804 27858
rect 6748 27188 6804 27806
rect 6748 27122 6804 27132
rect 6860 25732 6916 30158
rect 6860 25666 6916 25676
rect 6972 26516 7028 38612
rect 7420 38162 7476 38892
rect 7420 38110 7422 38162
rect 7474 38110 7476 38162
rect 7420 38098 7476 38110
rect 7532 38050 7588 39564
rect 7756 39060 7812 39788
rect 7756 38834 7812 39004
rect 7756 38782 7758 38834
rect 7810 38782 7812 38834
rect 7756 38770 7812 38782
rect 7868 39788 8036 39844
rect 8092 40180 8148 40190
rect 8092 40068 8148 40124
rect 8316 40068 8372 42588
rect 8428 40404 8484 40414
rect 8540 40404 8596 43708
rect 8764 42756 8820 42766
rect 8764 42662 8820 42700
rect 8876 42644 8932 45724
rect 8988 42980 9044 46844
rect 9100 46788 9156 46798
rect 9212 46788 9268 47292
rect 9156 46732 9268 46788
rect 9100 46722 9156 46732
rect 9884 46004 9940 46014
rect 9884 45910 9940 45948
rect 9548 45892 9604 45902
rect 9324 45780 9380 45790
rect 9324 45686 9380 45724
rect 8988 42924 9156 42980
rect 8932 42588 9044 42644
rect 8876 42550 8932 42588
rect 8876 42196 8932 42206
rect 8876 42102 8932 42140
rect 8988 42082 9044 42588
rect 8988 42030 8990 42082
rect 9042 42030 9044 42082
rect 8988 42018 9044 42030
rect 9100 41188 9156 42924
rect 8428 40402 8596 40404
rect 8428 40350 8430 40402
rect 8482 40350 8596 40402
rect 8428 40348 8596 40350
rect 8764 41186 9156 41188
rect 8764 41134 9102 41186
rect 9154 41134 9156 41186
rect 8764 41132 9156 41134
rect 8764 40516 8820 41132
rect 9100 41122 9156 41132
rect 9324 42756 9380 42766
rect 9324 41186 9380 42700
rect 9324 41134 9326 41186
rect 9378 41134 9380 41186
rect 9324 41122 9380 41134
rect 9436 41860 9492 41870
rect 8428 40338 8484 40348
rect 8764 40290 8820 40460
rect 8764 40238 8766 40290
rect 8818 40238 8820 40290
rect 8764 40226 8820 40238
rect 9100 40402 9156 40414
rect 9100 40350 9102 40402
rect 9154 40350 9156 40402
rect 8092 40012 8372 40068
rect 7532 37998 7534 38050
rect 7586 37998 7588 38050
rect 7532 37986 7588 37998
rect 7644 38610 7700 38622
rect 7644 38558 7646 38610
rect 7698 38558 7700 38610
rect 7084 37828 7140 37838
rect 7084 36594 7140 37772
rect 7644 37268 7700 38558
rect 7756 37268 7812 37278
rect 7644 37266 7812 37268
rect 7644 37214 7758 37266
rect 7810 37214 7812 37266
rect 7644 37212 7812 37214
rect 7420 37156 7476 37166
rect 7420 37062 7476 37100
rect 7084 36542 7086 36594
rect 7138 36542 7140 36594
rect 7084 36530 7140 36542
rect 7644 35922 7700 37212
rect 7756 37202 7812 37212
rect 7868 36596 7924 39788
rect 8092 39730 8148 40012
rect 8092 39678 8094 39730
rect 8146 39678 8148 39730
rect 8092 39666 8148 39678
rect 8204 39844 8260 39854
rect 7980 39620 8036 39630
rect 7980 38834 8036 39564
rect 8204 39506 8260 39788
rect 8204 39454 8206 39506
rect 8258 39454 8260 39506
rect 8204 39442 8260 39454
rect 8316 39732 8372 39742
rect 7980 38782 7982 38834
rect 8034 38782 8036 38834
rect 7980 38770 8036 38782
rect 8092 38724 8148 38762
rect 8092 38658 8148 38668
rect 8204 38052 8260 38062
rect 8204 37490 8260 37996
rect 8204 37438 8206 37490
rect 8258 37438 8260 37490
rect 8204 37426 8260 37438
rect 8316 36820 8372 39676
rect 8652 38724 8708 38762
rect 8652 38658 8708 38668
rect 8988 37380 9044 37390
rect 8652 37268 8708 37278
rect 8540 37266 8708 37268
rect 8540 37214 8654 37266
rect 8706 37214 8708 37266
rect 8540 37212 8708 37214
rect 8204 36764 8372 36820
rect 8428 37156 8484 37166
rect 7980 36596 8036 36606
rect 7868 36594 8148 36596
rect 7868 36542 7982 36594
rect 8034 36542 8148 36594
rect 7868 36540 8148 36542
rect 7980 36530 8036 36540
rect 7644 35870 7646 35922
rect 7698 35870 7700 35922
rect 7644 35858 7700 35870
rect 7756 36148 7812 36158
rect 7644 34802 7700 34814
rect 7644 34750 7646 34802
rect 7698 34750 7700 34802
rect 7084 34020 7140 34030
rect 7308 34020 7364 34030
rect 7532 34020 7588 34030
rect 7084 34018 7532 34020
rect 7084 33966 7086 34018
rect 7138 33966 7310 34018
rect 7362 33966 7532 34018
rect 7084 33964 7532 33966
rect 7084 33954 7140 33964
rect 7308 33954 7364 33964
rect 7532 33954 7588 33964
rect 7084 33236 7140 33246
rect 7084 32004 7140 33180
rect 7420 33234 7476 33246
rect 7420 33182 7422 33234
rect 7474 33182 7476 33234
rect 7308 32564 7364 32574
rect 7308 32470 7364 32508
rect 7084 29652 7140 31948
rect 7420 31332 7476 33182
rect 7644 33012 7700 34750
rect 7756 33458 7812 36092
rect 8092 34916 8148 36540
rect 8204 36594 8260 36764
rect 8428 36708 8484 37100
rect 8204 36542 8206 36594
rect 8258 36542 8260 36594
rect 8204 36530 8260 36542
rect 8316 36652 8484 36708
rect 8204 35586 8260 35598
rect 8204 35534 8206 35586
rect 8258 35534 8260 35586
rect 8204 35364 8260 35534
rect 8204 35298 8260 35308
rect 8316 35252 8372 36652
rect 8540 35700 8596 37212
rect 8652 37202 8708 37212
rect 8764 37266 8820 37278
rect 8764 37214 8766 37266
rect 8818 37214 8820 37266
rect 8764 37044 8820 37214
rect 8988 37266 9044 37324
rect 8988 37214 8990 37266
rect 9042 37214 9044 37266
rect 8988 37202 9044 37214
rect 8988 37044 9044 37054
rect 8764 36988 8988 37044
rect 8988 36978 9044 36988
rect 8652 36482 8708 36494
rect 8652 36430 8654 36482
rect 8706 36430 8708 36482
rect 8652 36260 8708 36430
rect 8988 36260 9044 36270
rect 8652 36258 9044 36260
rect 8652 36206 8990 36258
rect 9042 36206 9044 36258
rect 8652 36204 9044 36206
rect 8988 35812 9044 36204
rect 8988 35746 9044 35756
rect 8540 35634 8596 35644
rect 8316 35196 8596 35252
rect 7868 34914 8148 34916
rect 7868 34862 8094 34914
rect 8146 34862 8148 34914
rect 7868 34860 8148 34862
rect 7868 34692 7924 34860
rect 8092 34850 8148 34860
rect 7868 34354 7924 34636
rect 7868 34302 7870 34354
rect 7922 34302 7924 34354
rect 7868 34290 7924 34302
rect 8092 34468 8148 34478
rect 7756 33406 7758 33458
rect 7810 33406 7812 33458
rect 7756 33394 7812 33406
rect 7644 32946 7700 32956
rect 7420 31266 7476 31276
rect 7532 31220 7588 31230
rect 7532 31126 7588 31164
rect 7980 30324 8036 30334
rect 7868 30210 7924 30222
rect 7868 30158 7870 30210
rect 7922 30158 7924 30210
rect 7532 30098 7588 30110
rect 7532 30046 7534 30098
rect 7586 30046 7588 30098
rect 7532 29764 7588 30046
rect 7756 29988 7812 29998
rect 7756 29894 7812 29932
rect 7868 29876 7924 30158
rect 7868 29810 7924 29820
rect 7532 29698 7588 29708
rect 7084 29650 7364 29652
rect 7084 29598 7086 29650
rect 7138 29598 7364 29650
rect 7084 29596 7364 29598
rect 7084 29586 7140 29596
rect 7308 29316 7364 29596
rect 7420 29540 7476 29550
rect 7420 29446 7476 29484
rect 7532 29426 7588 29438
rect 7980 29428 8036 30268
rect 7532 29374 7534 29426
rect 7586 29374 7588 29426
rect 7532 29316 7588 29374
rect 7308 29260 7588 29316
rect 7756 29426 8036 29428
rect 7756 29374 7982 29426
rect 8034 29374 8036 29426
rect 7756 29372 8036 29374
rect 7084 28530 7140 28542
rect 7084 28478 7086 28530
rect 7138 28478 7140 28530
rect 7084 28084 7140 28478
rect 7756 28532 7812 29372
rect 7980 29362 8036 29372
rect 7756 28466 7812 28476
rect 7980 28420 8036 28430
rect 7868 28418 8036 28420
rect 7868 28366 7982 28418
rect 8034 28366 8036 28418
rect 7868 28364 8036 28366
rect 7196 28084 7252 28094
rect 7084 28082 7252 28084
rect 7084 28030 7198 28082
rect 7250 28030 7252 28082
rect 7084 28028 7252 28030
rect 7196 28018 7252 28028
rect 7084 27860 7140 27870
rect 7084 27766 7140 27804
rect 7756 27860 7812 27870
rect 7756 27766 7812 27804
rect 7868 26628 7924 28364
rect 7980 28354 8036 28364
rect 7980 27970 8036 27982
rect 7980 27918 7982 27970
rect 8034 27918 8036 27970
rect 7980 27524 8036 27918
rect 7980 27458 8036 27468
rect 7868 26572 8036 26628
rect 7308 26516 7364 26526
rect 6972 26514 7364 26516
rect 6972 26462 6974 26514
rect 7026 26462 7310 26514
rect 7362 26462 7364 26514
rect 6972 26460 7364 26462
rect 6972 24948 7028 26460
rect 7308 26450 7364 26460
rect 7868 26404 7924 26414
rect 7868 26310 7924 26348
rect 7644 26292 7700 26302
rect 7308 25732 7364 25742
rect 7308 25638 7364 25676
rect 7084 25620 7140 25630
rect 7084 25526 7140 25564
rect 7532 25508 7588 25518
rect 7532 25414 7588 25452
rect 7644 25506 7700 26236
rect 7644 25454 7646 25506
rect 7698 25454 7700 25506
rect 7644 25442 7700 25454
rect 7756 25620 7812 25630
rect 7196 24948 7252 24958
rect 6972 24946 7252 24948
rect 6972 24894 6974 24946
rect 7026 24894 7198 24946
rect 7250 24894 7252 24946
rect 6972 24892 7252 24894
rect 6972 24882 7028 24892
rect 7196 24882 7252 24892
rect 7756 24722 7812 25564
rect 7868 25394 7924 25406
rect 7868 25342 7870 25394
rect 7922 25342 7924 25394
rect 7868 25284 7924 25342
rect 7868 25218 7924 25228
rect 7756 24670 7758 24722
rect 7810 24670 7812 24722
rect 7756 24658 7812 24670
rect 7980 21812 8036 26572
rect 7980 21746 8036 21756
rect 8092 20188 8148 34412
rect 8540 34356 8596 35196
rect 8540 34130 8596 34300
rect 8540 34078 8542 34130
rect 8594 34078 8596 34130
rect 8540 34066 8596 34078
rect 8652 34914 8708 34926
rect 8652 34862 8654 34914
rect 8706 34862 8708 34914
rect 8204 34020 8260 34030
rect 8316 34020 8372 34030
rect 8260 34018 8372 34020
rect 8260 33966 8318 34018
rect 8370 33966 8372 34018
rect 8260 33964 8372 33966
rect 8204 25060 8260 33964
rect 8316 33954 8372 33964
rect 8652 33348 8708 34862
rect 8652 33282 8708 33292
rect 8876 33906 8932 33918
rect 8876 33854 8878 33906
rect 8930 33854 8932 33906
rect 8428 33234 8484 33246
rect 8428 33182 8430 33234
rect 8482 33182 8484 33234
rect 8428 31668 8484 33182
rect 8876 32900 8932 33854
rect 8876 32834 8932 32844
rect 9100 32788 9156 40350
rect 9436 40292 9492 41804
rect 9548 41300 9604 45836
rect 10108 44100 10164 49196
rect 10220 49532 10556 49588
rect 10220 49138 10276 49532
rect 10220 49086 10222 49138
rect 10274 49086 10276 49138
rect 10220 49074 10276 49086
rect 10220 48356 10276 48366
rect 10220 48130 10276 48300
rect 10220 48078 10222 48130
rect 10274 48078 10276 48130
rect 10220 45892 10276 48078
rect 10332 46900 10388 46910
rect 10332 46786 10388 46844
rect 10332 46734 10334 46786
rect 10386 46734 10388 46786
rect 10332 46722 10388 46734
rect 10444 46676 10500 49532
rect 10556 49522 10612 49532
rect 10668 48804 10724 49756
rect 11228 49588 11284 49598
rect 11228 49494 11284 49532
rect 11116 49252 11172 49262
rect 11116 49158 11172 49196
rect 11340 49138 11396 49756
rect 11340 49086 11342 49138
rect 11394 49086 11396 49138
rect 11340 49074 11396 49086
rect 11452 49810 11844 49812
rect 11452 49758 11566 49810
rect 11618 49758 11844 49810
rect 11452 49756 11844 49758
rect 11452 49026 11508 49756
rect 11564 49746 11620 49756
rect 11788 49140 11844 49756
rect 12236 49810 12292 49980
rect 12572 49970 12628 49980
rect 12236 49758 12238 49810
rect 12290 49758 12292 49810
rect 12236 49746 12292 49758
rect 12908 49810 12964 50372
rect 12908 49758 12910 49810
rect 12962 49758 12964 49810
rect 11900 49588 11956 49598
rect 11900 49586 12068 49588
rect 11900 49534 11902 49586
rect 11954 49534 12068 49586
rect 11900 49532 12068 49534
rect 11900 49522 11956 49532
rect 11900 49140 11956 49150
rect 11788 49138 11956 49140
rect 11788 49086 11902 49138
rect 11954 49086 11956 49138
rect 11788 49084 11956 49086
rect 11900 49074 11956 49084
rect 11452 48974 11454 49026
rect 11506 48974 11508 49026
rect 11452 48962 11508 48974
rect 10668 48738 10724 48748
rect 11340 48804 11396 48814
rect 10780 48354 10836 48366
rect 10780 48302 10782 48354
rect 10834 48302 10836 48354
rect 10556 48244 10612 48254
rect 10556 48150 10612 48188
rect 10780 47460 10836 48302
rect 11340 48242 11396 48748
rect 11452 48356 11508 48366
rect 11508 48300 11732 48356
rect 11452 48290 11508 48300
rect 11340 48190 11342 48242
rect 11394 48190 11396 48242
rect 11340 48020 11396 48190
rect 11676 48244 11732 48300
rect 11788 48244 11844 48254
rect 11676 48242 11844 48244
rect 11676 48190 11790 48242
rect 11842 48190 11844 48242
rect 11676 48188 11844 48190
rect 11788 48178 11844 48188
rect 11676 48020 11732 48030
rect 11340 47964 11508 48020
rect 11340 47796 11396 47806
rect 10836 47404 11284 47460
rect 10780 47366 10836 47404
rect 10444 46674 11172 46676
rect 10444 46622 10446 46674
rect 10498 46622 11172 46674
rect 10444 46620 11172 46622
rect 10444 46610 10500 46620
rect 11004 46004 11060 46014
rect 10332 45892 10388 45902
rect 10220 45890 10388 45892
rect 10220 45838 10334 45890
rect 10386 45838 10388 45890
rect 10220 45836 10388 45838
rect 10220 45218 10276 45230
rect 10220 45166 10222 45218
rect 10274 45166 10276 45218
rect 10220 44884 10276 45166
rect 10332 44884 10388 45836
rect 10892 45892 10948 45902
rect 10892 45778 10948 45836
rect 10892 45726 10894 45778
rect 10946 45726 10948 45778
rect 10892 45714 10948 45726
rect 10444 45668 10500 45678
rect 10444 45574 10500 45612
rect 10780 45668 10836 45678
rect 10444 44884 10500 44894
rect 10220 44828 10444 44884
rect 10444 44818 10500 44828
rect 10556 44772 10612 44782
rect 10556 44660 10612 44716
rect 10220 44604 10612 44660
rect 10220 44322 10276 44604
rect 10220 44270 10222 44322
rect 10274 44270 10276 44322
rect 10220 44258 10276 44270
rect 10444 44324 10500 44334
rect 10444 44230 10500 44268
rect 10556 44210 10612 44222
rect 10556 44158 10558 44210
rect 10610 44158 10612 44210
rect 10556 44100 10612 44158
rect 10108 44044 10276 44100
rect 9996 43988 10052 43998
rect 9884 43932 9996 43988
rect 9548 41234 9604 41244
rect 9660 43314 9716 43326
rect 9660 43262 9662 43314
rect 9714 43262 9716 43314
rect 9660 42308 9716 43262
rect 9772 43314 9828 43326
rect 9772 43262 9774 43314
rect 9826 43262 9828 43314
rect 9772 42756 9828 43262
rect 9884 43204 9940 43932
rect 9996 43922 10052 43932
rect 10108 43540 10164 43550
rect 10108 43446 10164 43484
rect 9996 43428 10052 43438
rect 9996 43334 10052 43372
rect 9884 43148 10052 43204
rect 9772 42690 9828 42700
rect 9212 40236 9492 40292
rect 9548 41076 9604 41086
rect 9548 40962 9604 41020
rect 9548 40910 9550 40962
rect 9602 40910 9604 40962
rect 9212 38276 9268 40236
rect 9548 38668 9604 40910
rect 9660 40514 9716 42252
rect 9660 40462 9662 40514
rect 9714 40462 9716 40514
rect 9660 40450 9716 40462
rect 9884 41300 9940 41310
rect 9884 40516 9940 41244
rect 9884 40402 9940 40460
rect 9884 40350 9886 40402
rect 9938 40350 9940 40402
rect 9884 40338 9940 40350
rect 9436 38612 9492 38622
rect 9548 38612 9716 38668
rect 9212 38210 9268 38220
rect 9324 38556 9436 38612
rect 9212 38052 9268 38062
rect 9324 38052 9380 38556
rect 9436 38546 9492 38556
rect 9548 38052 9604 38062
rect 9212 38050 9380 38052
rect 9212 37998 9214 38050
rect 9266 37998 9380 38050
rect 9212 37996 9380 37998
rect 9436 38050 9604 38052
rect 9436 37998 9550 38050
rect 9602 37998 9604 38050
rect 9436 37996 9604 37998
rect 9212 37380 9268 37996
rect 9212 37314 9268 37324
rect 9212 33460 9268 33470
rect 9212 33346 9268 33404
rect 9212 33294 9214 33346
rect 9266 33294 9268 33346
rect 9212 33282 9268 33294
rect 9100 32732 9268 32788
rect 8988 32564 9044 32574
rect 8988 32562 9156 32564
rect 8988 32510 8990 32562
rect 9042 32510 9156 32562
rect 8988 32508 9156 32510
rect 8988 32498 9044 32508
rect 8540 32450 8596 32462
rect 8540 32398 8542 32450
rect 8594 32398 8596 32450
rect 8540 31780 8596 32398
rect 9100 31892 9156 32508
rect 9100 31826 9156 31836
rect 8988 31780 9044 31790
rect 8540 31778 9044 31780
rect 8540 31726 8990 31778
rect 9042 31726 9044 31778
rect 8540 31724 9044 31726
rect 8428 31602 8484 31612
rect 8988 30996 9044 31724
rect 9100 31444 9156 31454
rect 9100 31218 9156 31388
rect 9100 31166 9102 31218
rect 9154 31166 9156 31218
rect 9100 31154 9156 31166
rect 8652 30882 8708 30894
rect 8652 30830 8654 30882
rect 8706 30830 8708 30882
rect 8652 30770 8708 30830
rect 8652 30718 8654 30770
rect 8706 30718 8708 30770
rect 8652 30706 8708 30718
rect 8652 30210 8708 30222
rect 8652 30158 8654 30210
rect 8706 30158 8708 30210
rect 8652 30100 8708 30158
rect 8540 29316 8596 29326
rect 8540 28308 8596 29260
rect 8652 28644 8708 30044
rect 8652 28578 8708 28588
rect 8876 29426 8932 29438
rect 8876 29374 8878 29426
rect 8930 29374 8932 29426
rect 8876 28644 8932 29374
rect 8876 28578 8932 28588
rect 8540 28082 8596 28252
rect 8764 28420 8820 28430
rect 8540 28030 8542 28082
rect 8594 28030 8596 28082
rect 8540 28018 8596 28030
rect 8652 28084 8708 28122
rect 8652 28018 8708 28028
rect 8764 28082 8820 28364
rect 8764 28030 8766 28082
rect 8818 28030 8820 28082
rect 8764 28018 8820 28030
rect 8876 28308 8932 28318
rect 8428 27860 8484 27870
rect 8428 27858 8596 27860
rect 8428 27806 8430 27858
rect 8482 27806 8596 27858
rect 8428 27804 8596 27806
rect 8428 27794 8484 27804
rect 8540 27524 8596 27804
rect 8540 27458 8596 27468
rect 8652 27748 8708 27758
rect 8652 25618 8708 27692
rect 8876 27186 8932 28252
rect 8988 27970 9044 30940
rect 9100 30770 9156 30782
rect 9100 30718 9102 30770
rect 9154 30718 9156 30770
rect 9100 30210 9156 30718
rect 9100 30158 9102 30210
rect 9154 30158 9156 30210
rect 9100 28868 9156 30158
rect 9212 29988 9268 32732
rect 9324 31778 9380 31790
rect 9324 31726 9326 31778
rect 9378 31726 9380 31778
rect 9324 30100 9380 31726
rect 9436 31444 9492 37996
rect 9548 37986 9604 37996
rect 9660 37828 9716 38612
rect 9548 37772 9716 37828
rect 9772 38276 9828 38286
rect 9548 31892 9604 37772
rect 9772 37378 9828 38220
rect 9996 38050 10052 43148
rect 10220 39620 10276 44044
rect 10444 44044 10612 44100
rect 10444 43092 10500 44044
rect 10444 43026 10500 43036
rect 10556 43876 10612 43886
rect 10332 42532 10388 42542
rect 10332 42438 10388 42476
rect 10556 42084 10612 43820
rect 10780 42756 10836 45612
rect 11004 44548 11060 45948
rect 11116 45106 11172 46620
rect 11228 45780 11284 47404
rect 11340 46786 11396 47740
rect 11452 46900 11508 47964
rect 11676 47926 11732 47964
rect 11788 47572 11844 47582
rect 11452 46844 11620 46900
rect 11340 46734 11342 46786
rect 11394 46734 11396 46786
rect 11340 46722 11396 46734
rect 11452 46676 11508 46686
rect 11452 46582 11508 46620
rect 11340 45780 11396 45790
rect 11228 45724 11340 45780
rect 11116 45054 11118 45106
rect 11170 45054 11172 45106
rect 11116 44772 11172 45054
rect 11116 44706 11172 44716
rect 11228 44884 11284 44894
rect 11004 44492 11172 44548
rect 11004 44324 11060 44334
rect 11004 44230 11060 44268
rect 11004 43652 11060 43662
rect 11004 43558 11060 43596
rect 10780 42662 10836 42700
rect 10892 42644 10948 42654
rect 10556 42028 10724 42084
rect 10332 41186 10388 41198
rect 10332 41134 10334 41186
rect 10386 41134 10388 41186
rect 10332 39844 10388 41134
rect 10332 39778 10388 39788
rect 10556 40740 10612 40750
rect 10556 40404 10612 40684
rect 10332 39620 10388 39630
rect 10220 39564 10332 39620
rect 10332 39554 10388 39564
rect 10556 39618 10612 40348
rect 10556 39566 10558 39618
rect 10610 39566 10612 39618
rect 10556 39554 10612 39566
rect 10556 39284 10612 39294
rect 10556 39060 10612 39228
rect 10332 39004 10612 39060
rect 10332 38668 10388 39004
rect 10668 38668 10724 42028
rect 10892 41186 10948 42588
rect 10892 41134 10894 41186
rect 10946 41134 10948 41186
rect 10892 41122 10948 41134
rect 11116 42082 11172 44492
rect 11228 44322 11284 44828
rect 11228 44270 11230 44322
rect 11282 44270 11284 44322
rect 11228 44258 11284 44270
rect 11340 44324 11396 45724
rect 11452 45668 11508 45678
rect 11564 45668 11620 46844
rect 11508 45612 11620 45668
rect 11452 45602 11508 45612
rect 11452 45164 11732 45220
rect 11452 45106 11508 45164
rect 11452 45054 11454 45106
rect 11506 45054 11508 45106
rect 11452 45042 11508 45054
rect 11564 44994 11620 45006
rect 11564 44942 11566 44994
rect 11618 44942 11620 44994
rect 11452 44324 11508 44334
rect 11340 44322 11508 44324
rect 11340 44270 11454 44322
rect 11506 44270 11508 44322
rect 11340 44268 11508 44270
rect 11452 44258 11508 44268
rect 11340 43764 11396 43774
rect 11340 43426 11396 43708
rect 11340 43374 11342 43426
rect 11394 43374 11396 43426
rect 11340 43362 11396 43374
rect 11452 43316 11508 43326
rect 11452 43222 11508 43260
rect 11116 42030 11118 42082
rect 11170 42030 11172 42082
rect 11116 39732 11172 42030
rect 11340 43092 11396 43102
rect 11340 42420 11396 43036
rect 11340 40404 11396 42364
rect 11452 41970 11508 41982
rect 11452 41918 11454 41970
rect 11506 41918 11508 41970
rect 11452 40740 11508 41918
rect 11452 40674 11508 40684
rect 11228 40348 11396 40404
rect 11452 40404 11508 40414
rect 11228 40180 11284 40348
rect 11452 40310 11508 40348
rect 11564 40180 11620 44942
rect 11676 43764 11732 45164
rect 11676 41972 11732 43708
rect 11788 43428 11844 47516
rect 12012 46004 12068 49532
rect 12796 48916 12852 48926
rect 12460 48804 12516 48814
rect 12460 48710 12516 48748
rect 12124 47572 12180 47582
rect 12180 47516 12292 47572
rect 12124 47506 12180 47516
rect 12236 47346 12292 47516
rect 12796 47458 12852 48860
rect 12908 48804 12964 49758
rect 12908 48738 12964 48748
rect 12796 47406 12798 47458
rect 12850 47406 12852 47458
rect 12796 47394 12852 47406
rect 12236 47294 12238 47346
rect 12290 47294 12292 47346
rect 12236 47282 12292 47294
rect 12684 47234 12740 47246
rect 12684 47182 12686 47234
rect 12738 47182 12740 47234
rect 12012 45938 12068 45948
rect 12572 46564 12628 46574
rect 12124 45890 12180 45902
rect 12124 45838 12126 45890
rect 12178 45838 12180 45890
rect 12124 45780 12180 45838
rect 12124 45714 12180 45724
rect 12236 44098 12292 44110
rect 12236 44046 12238 44098
rect 12290 44046 12292 44098
rect 11788 42644 11844 43372
rect 12124 43652 12180 43662
rect 11900 43316 11956 43326
rect 11956 43260 12068 43316
rect 11900 43250 11956 43260
rect 11900 42644 11956 42654
rect 11844 42642 11956 42644
rect 11844 42590 11902 42642
rect 11954 42590 11956 42642
rect 11844 42588 11956 42590
rect 11788 42550 11844 42588
rect 11900 42578 11956 42588
rect 11676 41916 11956 41972
rect 11900 41186 11956 41916
rect 11900 41134 11902 41186
rect 11954 41134 11956 41186
rect 11900 41122 11956 41134
rect 12012 40964 12068 43260
rect 12124 42082 12180 43596
rect 12236 42308 12292 44046
rect 12460 43428 12516 43438
rect 12460 43334 12516 43372
rect 12236 42242 12292 42252
rect 12124 42030 12126 42082
rect 12178 42030 12180 42082
rect 12124 41074 12180 42030
rect 12236 41970 12292 41982
rect 12236 41918 12238 41970
rect 12290 41918 12292 41970
rect 12236 41636 12292 41918
rect 12236 41580 12404 41636
rect 12124 41022 12126 41074
rect 12178 41022 12180 41074
rect 12124 41010 12180 41022
rect 11900 40908 12068 40964
rect 12236 40964 12292 40974
rect 11676 40516 11732 40526
rect 11676 40422 11732 40460
rect 11228 40124 11396 40180
rect 10892 39730 11172 39732
rect 10892 39678 11118 39730
rect 11170 39678 11172 39730
rect 10892 39676 11172 39678
rect 10780 39620 10836 39630
rect 10780 38836 10836 39564
rect 10780 38770 10836 38780
rect 10332 38612 10500 38668
rect 10668 38612 10836 38668
rect 9996 37998 9998 38050
rect 10050 37998 10052 38050
rect 9996 37986 10052 37998
rect 9772 37326 9774 37378
rect 9826 37326 9828 37378
rect 9772 37314 9828 37326
rect 9660 37266 9716 37278
rect 9660 37214 9662 37266
rect 9714 37214 9716 37266
rect 9660 37044 9716 37214
rect 9660 34580 9716 36988
rect 9884 37266 9940 37278
rect 9884 37214 9886 37266
rect 9938 37214 9940 37266
rect 9772 35698 9828 35710
rect 9772 35646 9774 35698
rect 9826 35646 9828 35698
rect 9772 35476 9828 35646
rect 9772 35410 9828 35420
rect 9884 35308 9940 37214
rect 10108 37268 10164 37278
rect 10108 37174 10164 37212
rect 10332 36260 10388 36270
rect 10108 35924 10164 35962
rect 10108 35858 10164 35868
rect 10332 35810 10388 36204
rect 10444 35922 10500 38612
rect 10556 38052 10612 38062
rect 10556 37490 10612 37996
rect 10668 37826 10724 37838
rect 10668 37774 10670 37826
rect 10722 37774 10724 37826
rect 10668 37716 10724 37774
rect 10668 37650 10724 37660
rect 10556 37438 10558 37490
rect 10610 37438 10612 37490
rect 10556 37426 10612 37438
rect 10556 36260 10612 36270
rect 10556 36166 10612 36204
rect 10444 35870 10446 35922
rect 10498 35870 10500 35922
rect 10444 35858 10500 35870
rect 10780 35812 10836 38612
rect 10892 37938 10948 39676
rect 11116 39666 11172 39676
rect 11004 39396 11060 39406
rect 11004 39302 11060 39340
rect 11228 39172 11284 39182
rect 11228 38276 11284 39116
rect 11228 38182 11284 38220
rect 10892 37886 10894 37938
rect 10946 37886 10948 37938
rect 10892 37874 10948 37886
rect 11340 37938 11396 40124
rect 11340 37886 11342 37938
rect 11394 37886 11396 37938
rect 11116 37826 11172 37838
rect 11116 37774 11118 37826
rect 11170 37774 11172 37826
rect 11116 37716 11172 37774
rect 11116 37044 11172 37660
rect 11116 36978 11172 36988
rect 10332 35758 10334 35810
rect 10386 35758 10388 35810
rect 10332 35746 10388 35758
rect 10668 35756 10836 35812
rect 11116 36260 11172 36270
rect 10444 35700 10500 35710
rect 10444 35588 10500 35644
rect 10332 35532 10500 35588
rect 10220 35308 10276 35318
rect 9884 35252 10052 35308
rect 9884 35028 9940 35038
rect 9884 34934 9940 34972
rect 9660 34514 9716 34524
rect 9660 34356 9716 34366
rect 9660 34130 9716 34300
rect 9660 34078 9662 34130
rect 9714 34078 9716 34130
rect 9660 34066 9716 34078
rect 9660 33460 9716 33470
rect 9660 33366 9716 33404
rect 9548 31826 9604 31836
rect 9660 32900 9716 32910
rect 9660 31778 9716 32844
rect 9660 31726 9662 31778
rect 9714 31726 9716 31778
rect 9660 31714 9716 31726
rect 9492 31388 9940 31444
rect 9436 31378 9492 31388
rect 9884 30210 9940 31388
rect 9884 30158 9886 30210
rect 9938 30158 9940 30210
rect 9660 30100 9716 30110
rect 9324 30098 9716 30100
rect 9324 30046 9662 30098
rect 9714 30046 9716 30098
rect 9324 30044 9716 30046
rect 9212 29932 9492 29988
rect 9100 28802 9156 28812
rect 8988 27918 8990 27970
rect 9042 27918 9044 27970
rect 8988 27906 9044 27918
rect 8876 27134 8878 27186
rect 8930 27134 8932 27186
rect 8876 27122 8932 27134
rect 8988 27748 9044 27758
rect 8652 25566 8654 25618
rect 8706 25566 8708 25618
rect 8652 25554 8708 25566
rect 8988 25506 9044 27692
rect 9212 27188 9268 27198
rect 9212 27094 9268 27132
rect 9100 27076 9156 27086
rect 9100 26982 9156 27020
rect 9324 26852 9380 26862
rect 9324 26758 9380 26796
rect 8988 25454 8990 25506
rect 9042 25454 9044 25506
rect 8988 25442 9044 25454
rect 9436 25506 9492 29932
rect 9660 29876 9716 30044
rect 9660 29810 9716 29820
rect 9772 29538 9828 29550
rect 9772 29486 9774 29538
rect 9826 29486 9828 29538
rect 9660 29428 9716 29438
rect 9660 29334 9716 29372
rect 9772 28084 9828 29486
rect 9772 28018 9828 28028
rect 9772 27074 9828 27086
rect 9772 27022 9774 27074
rect 9826 27022 9828 27074
rect 9772 26964 9828 27022
rect 9772 26898 9828 26908
rect 9548 26852 9604 26862
rect 9548 26290 9604 26796
rect 9660 26516 9716 26526
rect 9660 26422 9716 26460
rect 9772 26516 9828 26526
rect 9884 26516 9940 30158
rect 9996 29988 10052 35252
rect 10108 35252 10220 35308
rect 10108 34356 10164 35252
rect 10220 35242 10276 35252
rect 10108 34244 10164 34300
rect 10108 34188 10276 34244
rect 10108 34020 10164 34030
rect 10108 33122 10164 33964
rect 10108 33070 10110 33122
rect 10162 33070 10164 33122
rect 10108 32228 10164 33070
rect 10108 32162 10164 32172
rect 10108 30996 10164 31006
rect 10108 30902 10164 30940
rect 9996 29922 10052 29932
rect 10220 29652 10276 34188
rect 10108 29596 10276 29652
rect 10332 34130 10388 35532
rect 10556 35476 10612 35486
rect 10444 35420 10556 35476
rect 10444 34914 10500 35420
rect 10556 35410 10612 35420
rect 10444 34862 10446 34914
rect 10498 34862 10500 34914
rect 10444 34850 10500 34862
rect 10668 34468 10724 35756
rect 10332 34078 10334 34130
rect 10386 34078 10388 34130
rect 10108 27860 10164 29596
rect 10220 29428 10276 29438
rect 10332 29428 10388 34078
rect 10444 34412 10724 34468
rect 10780 35586 10836 35598
rect 10780 35534 10782 35586
rect 10834 35534 10836 35586
rect 10780 35476 10836 35534
rect 11116 35476 11172 36204
rect 10444 33460 10500 34412
rect 10556 34244 10612 34254
rect 10556 34150 10612 34188
rect 10668 34130 10724 34142
rect 10668 34078 10670 34130
rect 10722 34078 10724 34130
rect 10668 34020 10724 34078
rect 10668 33954 10724 33964
rect 10780 33684 10836 35420
rect 10892 35420 11172 35476
rect 10892 34914 10948 35420
rect 10892 34862 10894 34914
rect 10946 34862 10948 34914
rect 10892 34850 10948 34862
rect 11004 34802 11060 34814
rect 11004 34750 11006 34802
rect 11058 34750 11060 34802
rect 10780 33628 10948 33684
rect 10444 33394 10500 33404
rect 10780 33460 10836 33470
rect 10668 33124 10724 33134
rect 10444 32564 10500 32574
rect 10444 29988 10500 32508
rect 10668 32450 10724 33068
rect 10668 32398 10670 32450
rect 10722 32398 10724 32450
rect 10668 30212 10724 32398
rect 10780 32338 10836 33404
rect 10892 32676 10948 33628
rect 10892 32610 10948 32620
rect 10780 32286 10782 32338
rect 10834 32286 10836 32338
rect 10780 32274 10836 32286
rect 11004 32340 11060 34750
rect 11116 34804 11172 34814
rect 11116 34802 11284 34804
rect 11116 34750 11118 34802
rect 11170 34750 11284 34802
rect 11116 34748 11284 34750
rect 11116 34738 11172 34748
rect 11116 34244 11172 34254
rect 11116 34018 11172 34188
rect 11116 33966 11118 34018
rect 11170 33966 11172 34018
rect 11116 33796 11172 33966
rect 11116 33730 11172 33740
rect 11004 32274 11060 32284
rect 11004 31778 11060 31790
rect 11004 31726 11006 31778
rect 11058 31726 11060 31778
rect 10892 31668 10948 31678
rect 10892 31218 10948 31612
rect 10892 31166 10894 31218
rect 10946 31166 10948 31218
rect 10892 31154 10948 31166
rect 11004 31444 11060 31726
rect 11004 30994 11060 31388
rect 11004 30942 11006 30994
rect 11058 30942 11060 30994
rect 11004 30930 11060 30942
rect 11228 30436 11284 34748
rect 11340 34692 11396 37886
rect 11340 34626 11396 34636
rect 11452 40124 11620 40180
rect 11788 40292 11844 40302
rect 11452 30548 11508 40124
rect 11788 39058 11844 40236
rect 11900 40290 11956 40908
rect 11900 40238 11902 40290
rect 11954 40238 11956 40290
rect 11900 40226 11956 40238
rect 12124 40852 12180 40862
rect 11788 39006 11790 39058
rect 11842 39006 11844 39058
rect 11788 38668 11844 39006
rect 12124 38668 12180 40796
rect 12236 40626 12292 40908
rect 12236 40574 12238 40626
rect 12290 40574 12292 40626
rect 12236 40562 12292 40574
rect 12236 39620 12292 39630
rect 12348 39620 12404 41580
rect 12572 41298 12628 46508
rect 12684 43988 12740 47182
rect 12684 43764 12740 43932
rect 12684 43698 12740 43708
rect 12796 46788 12852 46798
rect 12796 43538 12852 46732
rect 13020 45220 13076 52334
rect 14588 52276 14644 54462
rect 15036 54514 15092 54526
rect 15036 54462 15038 54514
rect 15090 54462 15092 54514
rect 15036 53508 15092 54462
rect 15708 54516 15764 54526
rect 15932 54516 15988 54526
rect 16268 54516 16324 55356
rect 16380 55346 16436 55356
rect 16828 55300 16884 55310
rect 15708 54514 15876 54516
rect 15708 54462 15710 54514
rect 15762 54462 15876 54514
rect 15708 54460 15876 54462
rect 15708 54450 15764 54460
rect 15484 53508 15540 53518
rect 15036 53506 15540 53508
rect 15036 53454 15486 53506
rect 15538 53454 15540 53506
rect 15036 53452 15540 53454
rect 14588 52162 14644 52220
rect 14588 52110 14590 52162
rect 14642 52110 14644 52162
rect 14588 52098 14644 52110
rect 14812 52500 14868 52510
rect 14812 52162 14868 52444
rect 14812 52110 14814 52162
rect 14866 52110 14868 52162
rect 14812 52098 14868 52110
rect 13244 51940 13300 51950
rect 13244 51378 13300 51884
rect 14700 51938 14756 51950
rect 14700 51886 14702 51938
rect 14754 51886 14756 51938
rect 14700 51716 14756 51886
rect 13916 51660 14756 51716
rect 13916 51490 13972 51660
rect 15036 51604 15092 53452
rect 15484 53060 15540 53452
rect 15484 52994 15540 53004
rect 15372 52834 15428 52846
rect 15372 52782 15374 52834
rect 15426 52782 15428 52834
rect 15372 52500 15428 52782
rect 15372 52434 15428 52444
rect 15820 52276 15876 54460
rect 15932 54514 16324 54516
rect 15932 54462 15934 54514
rect 15986 54462 16324 54514
rect 15932 54460 16324 54462
rect 16380 54516 16436 54526
rect 16380 54514 16548 54516
rect 16380 54462 16382 54514
rect 16434 54462 16548 54514
rect 16380 54460 16548 54462
rect 15932 53284 15988 54460
rect 16380 54450 16436 54460
rect 16044 53844 16100 53854
rect 16044 53508 16100 53788
rect 16380 53508 16436 53518
rect 16044 53506 16436 53508
rect 16044 53454 16046 53506
rect 16098 53454 16382 53506
rect 16434 53454 16436 53506
rect 16044 53452 16436 53454
rect 16492 53508 16548 54460
rect 16716 53508 16772 53518
rect 16492 53506 16772 53508
rect 16492 53454 16718 53506
rect 16770 53454 16772 53506
rect 16492 53452 16772 53454
rect 16044 53442 16100 53452
rect 16380 53396 16436 53452
rect 16380 53340 16548 53396
rect 15932 53228 16100 53284
rect 15596 52220 15876 52276
rect 15596 52162 15652 52220
rect 15596 52110 15598 52162
rect 15650 52110 15652 52162
rect 15148 52050 15204 52062
rect 15148 51998 15150 52050
rect 15202 51998 15204 52050
rect 15148 51940 15204 51998
rect 15596 52052 15652 52110
rect 15596 51986 15652 51996
rect 15148 51874 15204 51884
rect 15708 51940 15764 51950
rect 15708 51846 15764 51884
rect 15820 51940 15876 51950
rect 15820 51938 15988 51940
rect 15820 51886 15822 51938
rect 15874 51886 15988 51938
rect 15820 51884 15988 51886
rect 15820 51874 15876 51884
rect 15036 51538 15092 51548
rect 13916 51438 13918 51490
rect 13970 51438 13972 51490
rect 13916 51426 13972 51438
rect 13244 51326 13246 51378
rect 13298 51326 13300 51378
rect 13244 50484 13300 51326
rect 15932 51268 15988 51884
rect 16044 51828 16100 53228
rect 16156 52948 16212 52958
rect 16156 52276 16212 52892
rect 16492 52724 16548 53340
rect 16492 52658 16548 52668
rect 16156 51940 16212 52220
rect 16268 52164 16324 52174
rect 16268 52070 16324 52108
rect 16492 52164 16548 52174
rect 16716 52164 16772 53452
rect 16548 52108 16772 52164
rect 16492 52098 16548 52108
rect 16828 52052 16884 55244
rect 17276 54514 17332 54526
rect 17276 54462 17278 54514
rect 17330 54462 17332 54514
rect 17276 52948 17332 54462
rect 17500 53396 17556 56140
rect 19180 56194 19236 56206
rect 19180 56142 19182 56194
rect 19234 56142 19236 56194
rect 18508 55412 18564 55422
rect 17724 55300 17780 55310
rect 17724 55206 17780 55244
rect 18396 55188 18452 55198
rect 17836 55186 18452 55188
rect 17836 55134 18398 55186
rect 18450 55134 18452 55186
rect 17836 55132 18452 55134
rect 17836 54852 17892 55132
rect 18396 55122 18452 55132
rect 17612 54796 17892 54852
rect 17612 54738 17668 54796
rect 17612 54686 17614 54738
rect 17666 54686 17668 54738
rect 17612 54674 17668 54686
rect 18508 54738 18564 55356
rect 18508 54686 18510 54738
rect 18562 54686 18564 54738
rect 18508 54674 18564 54686
rect 18732 54628 18788 54638
rect 18620 54626 18788 54628
rect 18620 54574 18734 54626
rect 18786 54574 18788 54626
rect 18620 54572 18788 54574
rect 17724 54514 17780 54526
rect 17724 54462 17726 54514
rect 17778 54462 17780 54514
rect 17724 53508 17780 54462
rect 17836 54516 17892 54526
rect 17836 54422 17892 54460
rect 18284 54514 18340 54526
rect 18284 54462 18286 54514
rect 18338 54462 18340 54514
rect 18172 53508 18228 53518
rect 17724 53452 18172 53508
rect 18172 53414 18228 53452
rect 17500 53340 18004 53396
rect 17276 52882 17332 52892
rect 17836 52274 17892 52286
rect 17836 52222 17838 52274
rect 17890 52222 17892 52274
rect 16604 51996 16884 52052
rect 17388 52052 17444 52062
rect 16156 51884 16548 51940
rect 16044 51772 16436 51828
rect 16044 51268 16100 51278
rect 15932 51266 16100 51268
rect 15932 51214 16046 51266
rect 16098 51214 16100 51266
rect 15932 51212 16100 51214
rect 15820 51156 15876 51166
rect 13244 50418 13300 50428
rect 15596 50596 15652 50606
rect 13132 50036 13188 50046
rect 13132 49942 13188 49980
rect 15484 49138 15540 49150
rect 15484 49086 15486 49138
rect 15538 49086 15540 49138
rect 15372 49028 15428 49038
rect 14476 48802 14532 48814
rect 14476 48750 14478 48802
rect 14530 48750 14532 48802
rect 14140 48244 14196 48254
rect 13804 48242 14196 48244
rect 13804 48190 14142 48242
rect 14194 48190 14196 48242
rect 13804 48188 14196 48190
rect 13468 48018 13524 48030
rect 13468 47966 13470 48018
rect 13522 47966 13524 48018
rect 13356 47684 13412 47694
rect 13132 47460 13188 47470
rect 13132 46788 13188 47404
rect 13356 46900 13412 47628
rect 13356 46806 13412 46844
rect 13468 46788 13524 47966
rect 13580 47458 13636 47470
rect 13580 47406 13582 47458
rect 13634 47406 13636 47458
rect 13580 47348 13636 47406
rect 13580 47282 13636 47292
rect 13804 47458 13860 48188
rect 14140 48178 14196 48188
rect 14364 48130 14420 48142
rect 14364 48078 14366 48130
rect 14418 48078 14420 48130
rect 13916 48020 13972 48030
rect 13916 47684 13972 47964
rect 13916 47628 14196 47684
rect 13804 47406 13806 47458
rect 13858 47406 13860 47458
rect 13804 47236 13860 47406
rect 14028 47460 14084 47470
rect 14028 47366 14084 47404
rect 13804 47180 14084 47236
rect 13468 46732 13636 46788
rect 13132 46694 13188 46732
rect 13580 46674 13636 46732
rect 13580 46622 13582 46674
rect 13634 46622 13636 46674
rect 13580 46564 13636 46622
rect 14028 46676 14084 47180
rect 14028 46610 14084 46620
rect 14140 46674 14196 47628
rect 14140 46622 14142 46674
rect 14194 46622 14196 46674
rect 14140 46610 14196 46622
rect 14252 47572 14308 47582
rect 13580 46508 13972 46564
rect 13916 45890 13972 46508
rect 13916 45838 13918 45890
rect 13970 45838 13972 45890
rect 13916 45826 13972 45838
rect 14252 45332 14308 47516
rect 14364 47460 14420 48078
rect 14476 48132 14532 48750
rect 14476 47684 14532 48076
rect 14476 47618 14532 47628
rect 14924 48802 14980 48814
rect 14924 48750 14926 48802
rect 14978 48750 14980 48802
rect 14812 47460 14868 47470
rect 14364 47404 14644 47460
rect 14588 47348 14644 47404
rect 14812 47366 14868 47404
rect 14700 47348 14756 47358
rect 14588 47292 14700 47348
rect 14476 47234 14532 47246
rect 14476 47182 14478 47234
rect 14530 47182 14532 47234
rect 14476 47124 14532 47182
rect 14476 47058 14532 47068
rect 14700 46674 14756 47292
rect 14700 46622 14702 46674
rect 14754 46622 14756 46674
rect 14476 46116 14532 46126
rect 14476 46002 14532 46060
rect 14700 46114 14756 46622
rect 14924 46676 14980 48750
rect 15372 48242 15428 48972
rect 15372 48190 15374 48242
rect 15426 48190 15428 48242
rect 15372 48178 15428 48190
rect 15260 48132 15316 48142
rect 15260 48038 15316 48076
rect 15372 47460 15428 47470
rect 15372 47366 15428 47404
rect 15484 47124 15540 49086
rect 15596 48018 15652 50540
rect 15820 49250 15876 51100
rect 15932 50706 15988 51212
rect 16044 51202 16100 51212
rect 15932 50654 15934 50706
rect 15986 50654 15988 50706
rect 15932 50642 15988 50654
rect 16044 50372 16100 50382
rect 16044 50370 16324 50372
rect 16044 50318 16046 50370
rect 16098 50318 16324 50370
rect 16044 50316 16324 50318
rect 16044 50306 16100 50316
rect 15820 49198 15822 49250
rect 15874 49198 15876 49250
rect 15820 49186 15876 49198
rect 16156 48804 16212 48814
rect 15932 48802 16212 48804
rect 15932 48750 16158 48802
rect 16210 48750 16212 48802
rect 15932 48748 16212 48750
rect 15596 47966 15598 48018
rect 15650 47966 15652 48018
rect 15596 47954 15652 47966
rect 15820 48020 15876 48030
rect 15484 47058 15540 47068
rect 15708 47458 15764 47470
rect 15708 47406 15710 47458
rect 15762 47406 15764 47458
rect 15036 46676 15092 46714
rect 14924 46620 15036 46676
rect 15036 46610 15092 46620
rect 15708 46562 15764 47406
rect 15708 46510 15710 46562
rect 15762 46510 15764 46562
rect 15036 46452 15092 46462
rect 14700 46062 14702 46114
rect 14754 46062 14756 46114
rect 14700 46050 14756 46062
rect 14924 46450 15092 46452
rect 14924 46398 15038 46450
rect 15090 46398 15092 46450
rect 14924 46396 15092 46398
rect 14476 45950 14478 46002
rect 14530 45950 14532 46002
rect 14476 45938 14532 45950
rect 13692 45276 14308 45332
rect 13020 45164 13300 45220
rect 12796 43486 12798 43538
rect 12850 43486 12852 43538
rect 12796 43474 12852 43486
rect 13020 44436 13076 44446
rect 12572 41246 12574 41298
rect 12626 41246 12628 41298
rect 12572 41234 12628 41246
rect 12684 43092 12740 43102
rect 12292 39564 12404 39620
rect 12236 39554 12292 39564
rect 12348 38836 12404 38846
rect 12348 38742 12404 38780
rect 11788 38612 11956 38668
rect 11788 38050 11844 38062
rect 11788 37998 11790 38050
rect 11842 37998 11844 38050
rect 11788 37380 11844 37998
rect 11900 38050 11956 38612
rect 11900 37998 11902 38050
rect 11954 37998 11956 38050
rect 11900 37986 11956 37998
rect 12012 38612 12180 38668
rect 11900 37380 11956 37390
rect 11788 37324 11900 37380
rect 11900 37266 11956 37324
rect 11900 37214 11902 37266
rect 11954 37214 11956 37266
rect 11900 37202 11956 37214
rect 12012 36148 12068 38612
rect 12124 38276 12180 38286
rect 12124 37828 12180 38220
rect 12236 38164 12292 38174
rect 12236 38070 12292 38108
rect 12348 38052 12404 38062
rect 12348 38050 12516 38052
rect 12348 37998 12350 38050
rect 12402 37998 12516 38050
rect 12348 37996 12516 37998
rect 12348 37986 12404 37996
rect 12124 37734 12180 37772
rect 12348 37828 12404 37838
rect 12460 37828 12516 37996
rect 12684 37828 12740 43036
rect 13020 42084 13076 44380
rect 13244 43762 13300 45164
rect 13692 44436 13748 45276
rect 13804 45108 13860 45118
rect 13860 45052 14308 45108
rect 13804 45014 13860 45052
rect 13804 44436 13860 44446
rect 13244 43710 13246 43762
rect 13298 43710 13300 43762
rect 13244 43698 13300 43710
rect 13580 44434 13860 44436
rect 13580 44382 13806 44434
rect 13858 44382 13860 44434
rect 13580 44380 13860 44382
rect 13132 43652 13188 43662
rect 13132 43558 13188 43596
rect 13468 43540 13524 43550
rect 13580 43540 13636 44380
rect 13804 44370 13860 44380
rect 14252 44322 14308 45052
rect 14364 44996 14420 45006
rect 14364 44994 14644 44996
rect 14364 44942 14366 44994
rect 14418 44942 14644 44994
rect 14364 44940 14644 44942
rect 14364 44930 14420 44940
rect 14252 44270 14254 44322
rect 14306 44270 14308 44322
rect 14252 44258 14308 44270
rect 14476 44548 14532 44558
rect 13468 43538 13636 43540
rect 13468 43486 13470 43538
rect 13522 43486 13636 43538
rect 13468 43484 13636 43486
rect 13916 43540 13972 43550
rect 13468 43474 13524 43484
rect 13916 43446 13972 43484
rect 14476 43426 14532 44492
rect 14476 43374 14478 43426
rect 14530 43374 14532 43426
rect 13468 43316 13524 43326
rect 13468 42754 13524 43260
rect 13916 42868 13972 42878
rect 13468 42702 13470 42754
rect 13522 42702 13524 42754
rect 13468 42690 13524 42702
rect 13692 42866 13972 42868
rect 13692 42814 13918 42866
rect 13970 42814 13972 42866
rect 13692 42812 13972 42814
rect 13020 42028 13188 42084
rect 13020 41858 13076 41870
rect 13020 41806 13022 41858
rect 13074 41806 13076 41858
rect 13020 41300 13076 41806
rect 13020 40626 13076 41244
rect 13020 40574 13022 40626
rect 13074 40574 13076 40626
rect 13020 40562 13076 40574
rect 12796 40402 12852 40414
rect 12796 40350 12798 40402
rect 12850 40350 12852 40402
rect 12796 39508 12852 40350
rect 12908 40292 12964 40302
rect 12908 40198 12964 40236
rect 12796 39442 12852 39452
rect 13132 39284 13188 42028
rect 13580 41076 13636 41086
rect 13580 40982 13636 41020
rect 13356 40740 13412 40750
rect 13356 40402 13412 40684
rect 13356 40350 13358 40402
rect 13410 40350 13412 40402
rect 13356 40338 13412 40350
rect 13132 39218 13188 39228
rect 13020 39060 13076 39070
rect 13020 38966 13076 39004
rect 12796 38834 12852 38846
rect 12796 38782 12798 38834
rect 12850 38782 12852 38834
rect 12796 38164 12852 38782
rect 13692 38668 13748 42812
rect 13916 42802 13972 42812
rect 13580 38612 13748 38668
rect 13804 42308 13860 42318
rect 13804 41410 13860 42252
rect 13804 41358 13806 41410
rect 13858 41358 13860 41410
rect 12796 38098 12852 38108
rect 13356 38500 13412 38510
rect 13356 38162 13412 38444
rect 13356 38110 13358 38162
rect 13410 38110 13412 38162
rect 13356 38098 13412 38110
rect 13020 37940 13076 37950
rect 12796 37828 12852 37838
rect 12460 37826 12852 37828
rect 12460 37774 12798 37826
rect 12850 37774 12852 37826
rect 12460 37772 12852 37774
rect 12124 37378 12180 37390
rect 12124 37326 12126 37378
rect 12178 37326 12180 37378
rect 12124 37044 12180 37326
rect 12124 36978 12180 36988
rect 12012 36082 12068 36092
rect 12012 35924 12068 35934
rect 12012 35830 12068 35868
rect 12012 35700 12068 35710
rect 11564 35588 11620 35598
rect 11564 35586 11732 35588
rect 11564 35534 11566 35586
rect 11618 35534 11732 35586
rect 11564 35532 11732 35534
rect 11564 35522 11620 35532
rect 11676 35252 11732 35532
rect 12012 35474 12068 35644
rect 12012 35422 12014 35474
rect 12066 35422 12068 35474
rect 12012 35410 12068 35422
rect 12124 35698 12180 35710
rect 12124 35646 12126 35698
rect 12178 35646 12180 35698
rect 11676 35196 11844 35252
rect 11564 35140 11620 35150
rect 11620 35084 11732 35140
rect 11564 35074 11620 35084
rect 11564 34804 11620 34814
rect 11564 34710 11620 34748
rect 11564 34356 11620 34366
rect 11676 34356 11732 35084
rect 11788 34692 11844 35196
rect 12012 34692 12068 34702
rect 11788 34690 12068 34692
rect 11788 34638 12014 34690
rect 12066 34638 12068 34690
rect 11788 34636 12068 34638
rect 12012 34468 12068 34636
rect 12012 34402 12068 34412
rect 11564 34354 11676 34356
rect 11564 34302 11566 34354
rect 11618 34302 11676 34354
rect 11564 34300 11676 34302
rect 11564 34290 11620 34300
rect 11676 34262 11732 34300
rect 12124 34132 12180 35646
rect 12236 35140 12292 35150
rect 12236 34914 12292 35084
rect 12348 35138 12404 37772
rect 12796 37716 12852 37772
rect 12908 37716 12964 37726
rect 12796 37660 12908 37716
rect 12908 37650 12964 37660
rect 12572 37492 12628 37502
rect 13020 37492 13076 37884
rect 13468 37938 13524 37950
rect 13468 37886 13470 37938
rect 13522 37886 13524 37938
rect 12572 37490 13076 37492
rect 12572 37438 12574 37490
rect 12626 37438 13022 37490
rect 13074 37438 13076 37490
rect 12572 37436 13076 37438
rect 12572 37380 12628 37436
rect 13020 37426 13076 37436
rect 13244 37716 13300 37726
rect 12572 37314 12628 37324
rect 12908 37268 12964 37278
rect 12908 36594 12964 37212
rect 12908 36542 12910 36594
rect 12962 36542 12964 36594
rect 12908 36484 12964 36542
rect 12572 36428 12908 36484
rect 12572 36260 12628 36428
rect 12908 36418 12964 36428
rect 12572 35922 12628 36204
rect 12572 35870 12574 35922
rect 12626 35870 12628 35922
rect 12572 35858 12628 35870
rect 13132 36148 13188 36158
rect 13020 35588 13076 35598
rect 12348 35086 12350 35138
rect 12402 35086 12404 35138
rect 12348 35074 12404 35086
rect 12908 35586 13076 35588
rect 12908 35534 13022 35586
rect 13074 35534 13076 35586
rect 12908 35532 13076 35534
rect 12236 34862 12238 34914
rect 12290 34862 12292 34914
rect 12236 34850 12292 34862
rect 12572 34916 12628 34926
rect 12572 34822 12628 34860
rect 12908 34692 12964 35532
rect 13020 35522 13076 35532
rect 12796 34690 12964 34692
rect 12796 34638 12910 34690
rect 12962 34638 12964 34690
rect 12796 34636 12964 34638
rect 12460 34132 12516 34142
rect 12796 34132 12852 34636
rect 12908 34626 12964 34636
rect 13020 34356 13076 34366
rect 13132 34356 13188 36092
rect 13020 34354 13188 34356
rect 13020 34302 13022 34354
rect 13074 34302 13188 34354
rect 13020 34300 13188 34302
rect 12124 34130 12852 34132
rect 12124 34078 12462 34130
rect 12514 34078 12852 34130
rect 12124 34076 12852 34078
rect 12908 34130 12964 34142
rect 12908 34078 12910 34130
rect 12962 34078 12964 34130
rect 12460 34066 12516 34076
rect 12012 34020 12068 34030
rect 11900 31666 11956 31678
rect 11900 31614 11902 31666
rect 11954 31614 11956 31666
rect 11452 30482 11508 30492
rect 11788 30994 11844 31006
rect 11788 30942 11790 30994
rect 11842 30942 11844 30994
rect 11228 30370 11284 30380
rect 11564 30436 11620 30446
rect 11564 30322 11620 30380
rect 11564 30270 11566 30322
rect 11618 30270 11620 30322
rect 11564 30258 11620 30270
rect 10668 30156 11172 30212
rect 10444 29922 10500 29932
rect 10668 29986 10724 29998
rect 10668 29934 10670 29986
rect 10722 29934 10724 29986
rect 10668 29876 10724 29934
rect 10668 29810 10724 29820
rect 10892 29988 10948 29998
rect 10220 29426 10388 29428
rect 10220 29374 10222 29426
rect 10274 29374 10388 29426
rect 10220 29372 10388 29374
rect 10668 29428 10724 29438
rect 10220 29362 10276 29372
rect 10220 29202 10276 29214
rect 10220 29150 10222 29202
rect 10274 29150 10276 29202
rect 10220 28642 10276 29150
rect 10668 28756 10724 29372
rect 10780 28756 10836 28766
rect 10668 28754 10836 28756
rect 10668 28702 10782 28754
rect 10834 28702 10836 28754
rect 10668 28700 10836 28702
rect 10780 28690 10836 28700
rect 10220 28590 10222 28642
rect 10274 28590 10276 28642
rect 10220 28578 10276 28590
rect 10556 28644 10612 28654
rect 10612 28588 10724 28644
rect 10556 28578 10612 28588
rect 10108 27794 10164 27804
rect 10332 28530 10388 28542
rect 10332 28478 10334 28530
rect 10386 28478 10388 28530
rect 9996 27748 10052 27758
rect 9996 27654 10052 27692
rect 10108 26964 10164 27002
rect 10108 26898 10164 26908
rect 9772 26514 9884 26516
rect 9772 26462 9774 26514
rect 9826 26462 9884 26514
rect 9772 26460 9884 26462
rect 9772 26450 9828 26460
rect 9884 26422 9940 26460
rect 10220 26404 10276 26414
rect 9548 26238 9550 26290
rect 9602 26238 9604 26290
rect 9548 25732 9604 26238
rect 9548 25666 9604 25676
rect 9660 26292 9716 26302
rect 9436 25454 9438 25506
rect 9490 25454 9492 25506
rect 9436 25442 9492 25454
rect 9660 25620 9716 26236
rect 10220 26290 10276 26348
rect 10220 26238 10222 26290
rect 10274 26238 10276 26290
rect 10220 26226 10276 26238
rect 9660 25506 9716 25564
rect 9660 25454 9662 25506
rect 9714 25454 9716 25506
rect 9660 25442 9716 25454
rect 10220 25508 10276 25518
rect 10220 25414 10276 25452
rect 9548 25396 9604 25406
rect 9548 25302 9604 25340
rect 8204 24994 8260 25004
rect 8316 25284 8372 25294
rect 8316 24946 8372 25228
rect 8316 24894 8318 24946
rect 8370 24894 8372 24946
rect 8316 24882 8372 24894
rect 9884 25282 9940 25294
rect 9884 25230 9886 25282
rect 9938 25230 9940 25282
rect 9884 24052 9940 25230
rect 9884 23986 9940 23996
rect 10332 23380 10388 28478
rect 10668 28420 10724 28588
rect 10780 28420 10836 28430
rect 10668 28418 10836 28420
rect 10668 28366 10782 28418
rect 10834 28366 10836 28418
rect 10668 28364 10836 28366
rect 10780 28354 10836 28364
rect 10892 28420 10948 29932
rect 11004 29428 11060 29438
rect 11004 29334 11060 29372
rect 10892 28326 10948 28364
rect 11116 28530 11172 30156
rect 11452 30210 11508 30222
rect 11452 30158 11454 30210
rect 11506 30158 11508 30210
rect 11452 30100 11508 30158
rect 11340 30044 11508 30100
rect 11676 30098 11732 30110
rect 11676 30046 11678 30098
rect 11730 30046 11732 30098
rect 11116 28478 11118 28530
rect 11170 28478 11172 28530
rect 10556 28084 10612 28094
rect 10556 27186 10612 28028
rect 11116 28084 11172 28478
rect 11116 28018 11172 28028
rect 11228 29986 11284 29998
rect 11228 29934 11230 29986
rect 11282 29934 11284 29986
rect 11228 29764 11284 29934
rect 10780 27860 10836 27870
rect 10780 27766 10836 27804
rect 10556 27134 10558 27186
rect 10610 27134 10612 27186
rect 10556 27076 10612 27134
rect 10556 27010 10612 27020
rect 10556 26516 10612 26526
rect 10556 26180 10612 26460
rect 10556 26114 10612 26124
rect 11004 26404 11060 26414
rect 11004 25956 11060 26348
rect 11228 26292 11284 29708
rect 11340 29652 11396 30044
rect 11564 29988 11620 29998
rect 11676 29988 11732 30046
rect 11788 30100 11844 30942
rect 11900 30324 11956 31614
rect 12012 31108 12068 33964
rect 12124 33124 12180 33134
rect 12460 33124 12516 33134
rect 12124 33122 12516 33124
rect 12124 33070 12126 33122
rect 12178 33070 12462 33122
rect 12514 33070 12516 33122
rect 12124 33068 12516 33070
rect 12124 33058 12180 33068
rect 12460 32340 12516 33068
rect 12460 32274 12516 32284
rect 12460 32116 12516 32126
rect 12012 31052 12292 31108
rect 12124 30884 12180 30894
rect 11900 30258 11956 30268
rect 12012 30828 12124 30884
rect 11788 30034 11844 30044
rect 11620 29932 11732 29988
rect 11900 29986 11956 29998
rect 11900 29934 11902 29986
rect 11954 29934 11956 29986
rect 11564 29922 11620 29932
rect 11900 29764 11956 29934
rect 11900 29698 11956 29708
rect 11340 29596 11620 29652
rect 11564 29540 11620 29596
rect 11788 29540 11844 29550
rect 12012 29540 12068 30828
rect 12124 30818 12180 30828
rect 12124 30100 12180 30110
rect 12124 30006 12180 30044
rect 11564 29484 11788 29540
rect 11788 29446 11844 29484
rect 11900 29484 12068 29540
rect 11900 29428 11956 29484
rect 11340 28868 11396 28878
rect 11340 28642 11396 28812
rect 11900 28754 11956 29372
rect 12124 29428 12180 29438
rect 12236 29428 12292 31052
rect 12460 29764 12516 32060
rect 12460 29698 12516 29708
rect 12572 31108 12628 31118
rect 12572 30098 12628 31052
rect 12684 30772 12740 34076
rect 12908 34020 12964 34078
rect 12908 33954 12964 33964
rect 13020 33460 13076 34300
rect 13244 34244 13300 37660
rect 13020 33394 13076 33404
rect 13132 34188 13300 34244
rect 13356 37044 13412 37054
rect 13020 33124 13076 33134
rect 13020 33030 13076 33068
rect 12796 32562 12852 32574
rect 12796 32510 12798 32562
rect 12850 32510 12852 32562
rect 12796 32340 12852 32510
rect 12796 31778 12852 32284
rect 13132 32564 13188 34188
rect 13132 32004 13188 32508
rect 13132 31938 13188 31948
rect 13244 33684 13300 33694
rect 12796 31726 12798 31778
rect 12850 31726 12852 31778
rect 12796 31714 12852 31726
rect 12908 31556 12964 31566
rect 12908 31462 12964 31500
rect 13132 31332 13188 31342
rect 13132 31218 13188 31276
rect 13132 31166 13134 31218
rect 13186 31166 13188 31218
rect 13132 31154 13188 31166
rect 13244 30996 13300 33628
rect 13356 32116 13412 36988
rect 13468 35700 13524 37886
rect 13580 37268 13636 38612
rect 13692 37828 13748 37838
rect 13692 37734 13748 37772
rect 13692 37268 13748 37278
rect 13580 37212 13692 37268
rect 13580 37044 13636 37054
rect 13580 35924 13636 36988
rect 13692 36148 13748 37212
rect 13804 36708 13860 41358
rect 14252 42196 14308 42206
rect 14252 41410 14308 42140
rect 14252 41358 14254 41410
rect 14306 41358 14308 41410
rect 14252 41346 14308 41358
rect 14028 41188 14084 41198
rect 14028 41094 14084 41132
rect 14140 41076 14196 41086
rect 14140 39620 14196 41020
rect 14364 40404 14420 40414
rect 14364 40310 14420 40348
rect 14476 40180 14532 43374
rect 14028 39564 14196 39620
rect 14364 40124 14532 40180
rect 14028 39060 14084 39564
rect 14140 39396 14196 39406
rect 14140 39394 14308 39396
rect 14140 39342 14142 39394
rect 14194 39342 14308 39394
rect 14140 39340 14308 39342
rect 14140 39330 14196 39340
rect 13916 38834 13972 38846
rect 13916 38782 13918 38834
rect 13970 38782 13972 38834
rect 13916 38276 13972 38782
rect 13916 38210 13972 38220
rect 14028 38050 14084 39004
rect 14252 39284 14308 39340
rect 14028 37998 14030 38050
rect 14082 37998 14084 38050
rect 14028 37986 14084 37998
rect 14140 38388 14196 38398
rect 13916 37828 13972 37838
rect 13916 37734 13972 37772
rect 13916 37604 13972 37614
rect 13916 36820 13972 37548
rect 14140 37268 14196 38332
rect 14252 37380 14308 39228
rect 14364 37604 14420 40124
rect 14476 39508 14532 39518
rect 14476 38834 14532 39452
rect 14476 38782 14478 38834
rect 14530 38782 14532 38834
rect 14476 38770 14532 38782
rect 14476 38276 14532 38286
rect 14476 37938 14532 38220
rect 14476 37886 14478 37938
rect 14530 37886 14532 37938
rect 14476 37874 14532 37886
rect 14364 37538 14420 37548
rect 14252 37324 14532 37380
rect 14028 37212 14196 37268
rect 14028 37044 14084 37212
rect 14028 36978 14084 36988
rect 13916 36764 14084 36820
rect 13804 36652 13972 36708
rect 13804 36484 13860 36494
rect 13804 36370 13860 36428
rect 13804 36318 13806 36370
rect 13858 36318 13860 36370
rect 13804 36306 13860 36318
rect 13692 36082 13748 36092
rect 13916 35924 13972 36652
rect 14028 36484 14084 36764
rect 14140 36708 14196 36718
rect 14140 36614 14196 36652
rect 14364 36484 14420 36494
rect 14028 36428 14308 36484
rect 13580 35868 13860 35924
rect 13468 35634 13524 35644
rect 13468 34916 13524 34926
rect 13468 32786 13524 34860
rect 13580 34692 13636 34702
rect 13580 34598 13636 34636
rect 13804 34690 13860 35868
rect 13916 35698 13972 35868
rect 13916 35646 13918 35698
rect 13970 35646 13972 35698
rect 13916 35634 13972 35646
rect 14028 36258 14084 36270
rect 14028 36206 14030 36258
rect 14082 36206 14084 36258
rect 13804 34638 13806 34690
rect 13858 34638 13860 34690
rect 13804 34626 13860 34638
rect 13916 34580 13972 34590
rect 13916 34354 13972 34524
rect 13916 34302 13918 34354
rect 13970 34302 13972 34354
rect 13916 34290 13972 34302
rect 14028 33684 14084 36206
rect 14028 33618 14084 33628
rect 14140 35476 14196 35486
rect 14140 33460 14196 35420
rect 14252 34468 14308 36428
rect 14364 36390 14420 36428
rect 14364 35586 14420 35598
rect 14364 35534 14366 35586
rect 14418 35534 14420 35586
rect 14364 34692 14420 35534
rect 14476 34916 14532 37324
rect 14476 34850 14532 34860
rect 14364 34626 14420 34636
rect 14252 34402 14308 34412
rect 14252 34242 14308 34254
rect 14252 34190 14254 34242
rect 14306 34190 14308 34242
rect 14252 33572 14308 34190
rect 14252 33506 14308 33516
rect 14364 34132 14420 34142
rect 14588 34132 14644 44940
rect 14812 44660 14868 44670
rect 14812 44434 14868 44604
rect 14812 44382 14814 44434
rect 14866 44382 14868 44434
rect 14812 44370 14868 44382
rect 14924 41412 14980 46396
rect 15036 46386 15092 46396
rect 15708 46452 15764 46510
rect 15708 46386 15764 46396
rect 15036 46114 15092 46126
rect 15036 46062 15038 46114
rect 15090 46062 15092 46114
rect 15036 46002 15092 46062
rect 15036 45950 15038 46002
rect 15090 45950 15092 46002
rect 15036 45938 15092 45950
rect 15820 46116 15876 47964
rect 15260 44322 15316 44334
rect 15260 44270 15262 44322
rect 15314 44270 15316 44322
rect 15260 43764 15316 44270
rect 15708 44322 15764 44334
rect 15708 44270 15710 44322
rect 15762 44270 15764 44322
rect 15708 43988 15764 44270
rect 15708 43922 15764 43932
rect 15260 43698 15316 43708
rect 15596 43764 15652 43774
rect 14924 41346 14980 41356
rect 15148 42644 15204 42654
rect 15036 41188 15092 41198
rect 14700 40962 14756 40974
rect 14700 40910 14702 40962
rect 14754 40910 14756 40962
rect 14700 40068 14756 40910
rect 15036 40962 15092 41132
rect 15036 40910 15038 40962
rect 15090 40910 15092 40962
rect 14700 40002 14756 40012
rect 14812 40292 14868 40302
rect 15036 40292 15092 40910
rect 14812 40290 15092 40292
rect 14812 40238 14814 40290
rect 14866 40238 15092 40290
rect 14812 40236 15092 40238
rect 14700 39508 14756 39518
rect 14700 39414 14756 39452
rect 14812 39396 14868 40236
rect 15036 40068 15092 40078
rect 15036 39618 15092 40012
rect 15036 39566 15038 39618
rect 15090 39566 15092 39618
rect 15036 39554 15092 39566
rect 14812 39330 14868 39340
rect 15148 39394 15204 42588
rect 15148 39342 15150 39394
rect 15202 39342 15204 39394
rect 15148 39330 15204 39342
rect 15260 40516 15316 40526
rect 15036 39172 15092 39182
rect 15036 39058 15092 39116
rect 15260 39060 15316 40460
rect 15372 40402 15428 40414
rect 15372 40350 15374 40402
rect 15426 40350 15428 40402
rect 15372 40068 15428 40350
rect 15372 40002 15428 40012
rect 15596 40404 15652 43708
rect 15708 41074 15764 41086
rect 15708 41022 15710 41074
rect 15762 41022 15764 41074
rect 15708 40852 15764 41022
rect 15708 40786 15764 40796
rect 15036 39006 15038 39058
rect 15090 39006 15092 39058
rect 15036 38994 15092 39006
rect 15148 39058 15316 39060
rect 15148 39006 15262 39058
rect 15314 39006 15316 39058
rect 15148 39004 15316 39006
rect 14812 38834 14868 38846
rect 14812 38782 14814 38834
rect 14866 38782 14868 38834
rect 14812 38388 14868 38782
rect 14812 38322 14868 38332
rect 15148 38162 15204 39004
rect 15260 38994 15316 39004
rect 15484 38836 15540 38846
rect 15484 38742 15540 38780
rect 15372 38612 15428 38622
rect 15372 38610 15540 38612
rect 15372 38558 15374 38610
rect 15426 38558 15540 38610
rect 15372 38556 15540 38558
rect 15372 38546 15428 38556
rect 15148 38110 15150 38162
rect 15202 38110 15204 38162
rect 15148 38098 15204 38110
rect 15036 38050 15092 38062
rect 15036 37998 15038 38050
rect 15090 37998 15092 38050
rect 15036 37940 15092 37998
rect 15036 37874 15092 37884
rect 15148 37380 15204 37390
rect 15148 37266 15204 37324
rect 15148 37214 15150 37266
rect 15202 37214 15204 37266
rect 15148 37202 15204 37214
rect 15372 37268 15428 37278
rect 15484 37268 15540 38556
rect 15596 38050 15652 40348
rect 15708 39844 15764 39854
rect 15708 38388 15764 39788
rect 15820 38388 15876 46060
rect 15932 40514 15988 48748
rect 16156 48738 16212 48748
rect 16044 48244 16100 48254
rect 16044 47458 16100 48188
rect 16156 48130 16212 48142
rect 16156 48078 16158 48130
rect 16210 48078 16212 48130
rect 16156 48018 16212 48078
rect 16156 47966 16158 48018
rect 16210 47966 16212 48018
rect 16156 47954 16212 47966
rect 16044 47406 16046 47458
rect 16098 47406 16100 47458
rect 16044 47394 16100 47406
rect 16156 47682 16212 47694
rect 16156 47630 16158 47682
rect 16210 47630 16212 47682
rect 16156 47460 16212 47630
rect 16044 47124 16100 47134
rect 16044 45890 16100 47068
rect 16156 46898 16212 47404
rect 16156 46846 16158 46898
rect 16210 46846 16212 46898
rect 16156 46834 16212 46846
rect 16044 45838 16046 45890
rect 16098 45838 16100 45890
rect 16044 45826 16100 45838
rect 16268 45778 16324 50316
rect 16380 48914 16436 51772
rect 16492 51602 16548 51884
rect 16492 51550 16494 51602
rect 16546 51550 16548 51602
rect 16492 51538 16548 51550
rect 16492 50708 16548 50718
rect 16604 50708 16660 51996
rect 17052 51604 17108 51614
rect 16828 51378 16884 51390
rect 16828 51326 16830 51378
rect 16882 51326 16884 51378
rect 16828 51156 16884 51326
rect 16828 51090 16884 51100
rect 16492 50706 16660 50708
rect 16492 50654 16494 50706
rect 16546 50654 16660 50706
rect 16492 50652 16660 50654
rect 16492 50484 16548 50652
rect 17052 50428 17108 51548
rect 17388 51602 17444 51996
rect 17388 51550 17390 51602
rect 17442 51550 17444 51602
rect 17388 51538 17444 51550
rect 17724 51378 17780 51390
rect 17724 51326 17726 51378
rect 17778 51326 17780 51378
rect 17724 51156 17780 51326
rect 17724 51090 17780 51100
rect 16492 50418 16548 50428
rect 16828 50372 17108 50428
rect 17612 50484 17668 50494
rect 16380 48862 16382 48914
rect 16434 48862 16436 48914
rect 16380 48850 16436 48862
rect 16492 48914 16548 48926
rect 16492 48862 16494 48914
rect 16546 48862 16548 48914
rect 16492 48244 16548 48862
rect 16828 48580 16884 50372
rect 17612 49922 17668 50428
rect 17612 49870 17614 49922
rect 17666 49870 17668 49922
rect 17612 49858 17668 49870
rect 17836 49924 17892 52222
rect 17948 50372 18004 53340
rect 18060 52948 18116 52958
rect 18060 52854 18116 52892
rect 18172 52836 18228 52846
rect 18172 52742 18228 52780
rect 18284 52612 18340 54462
rect 18396 54516 18452 54526
rect 18396 54422 18452 54460
rect 18172 52556 18340 52612
rect 18396 52946 18452 52958
rect 18396 52894 18398 52946
rect 18450 52894 18452 52946
rect 18060 52276 18116 52286
rect 18060 50428 18116 52220
rect 18172 52052 18228 52556
rect 18396 52500 18452 52894
rect 18396 52434 18452 52444
rect 18508 52946 18564 52958
rect 18508 52894 18510 52946
rect 18562 52894 18564 52946
rect 18508 52164 18564 52894
rect 18172 51602 18228 51996
rect 18172 51550 18174 51602
rect 18226 51550 18228 51602
rect 18172 51538 18228 51550
rect 18284 52108 18564 52164
rect 18620 52164 18676 54572
rect 18732 54562 18788 54572
rect 19068 52834 19124 52846
rect 19068 52782 19070 52834
rect 19122 52782 19124 52834
rect 19068 52500 19124 52782
rect 19068 52434 19124 52444
rect 19180 52276 19236 56142
rect 20860 56196 20916 56252
rect 23100 56420 23156 59200
rect 25340 56420 25396 59200
rect 27580 57204 27636 59200
rect 27580 57148 27972 57204
rect 23100 56364 23604 56420
rect 23100 56306 23156 56364
rect 23100 56254 23102 56306
rect 23154 56254 23156 56306
rect 23100 56242 23156 56254
rect 21084 56196 21140 56206
rect 21420 56196 21476 56206
rect 20860 56194 21140 56196
rect 20860 56142 21086 56194
rect 21138 56142 21140 56194
rect 20860 56140 21140 56142
rect 21084 56130 21140 56140
rect 21308 56194 21476 56196
rect 21308 56142 21422 56194
rect 21474 56142 21476 56194
rect 21308 56140 21476 56142
rect 20524 55412 20580 55422
rect 20524 55318 20580 55356
rect 19836 54908 20100 54918
rect 19892 54852 19940 54908
rect 19996 54852 20044 54908
rect 19836 54842 20100 54852
rect 21084 54514 21140 54526
rect 21084 54462 21086 54514
rect 21138 54462 21140 54514
rect 19836 53340 20100 53350
rect 19892 53284 19940 53340
rect 19996 53284 20044 53340
rect 19836 53274 20100 53284
rect 19180 52210 19236 52220
rect 19964 52836 20020 52846
rect 19964 52274 20020 52780
rect 19964 52222 19966 52274
rect 20018 52222 20020 52274
rect 19964 52210 20020 52222
rect 18284 51602 18340 52108
rect 18284 51550 18286 51602
rect 18338 51550 18340 51602
rect 18284 51538 18340 51550
rect 18620 51602 18676 52108
rect 20636 52164 20692 52174
rect 20636 52070 20692 52108
rect 21084 52164 21140 54462
rect 19836 51772 20100 51782
rect 19892 51716 19940 51772
rect 19996 51716 20044 51772
rect 19836 51706 20100 51716
rect 18620 51550 18622 51602
rect 18674 51550 18676 51602
rect 18620 51538 18676 51550
rect 18396 51378 18452 51390
rect 18396 51326 18398 51378
rect 18450 51326 18452 51378
rect 18172 50482 18228 50494
rect 18172 50430 18174 50482
rect 18226 50430 18228 50482
rect 18172 50428 18228 50430
rect 18060 50372 18228 50428
rect 17948 50306 18004 50316
rect 17836 49858 17892 49868
rect 18172 49252 18228 50372
rect 16604 48524 16884 48580
rect 16604 48466 16660 48524
rect 16604 48414 16606 48466
rect 16658 48414 16660 48466
rect 16604 48402 16660 48414
rect 16492 48178 16548 48188
rect 16380 48018 16436 48030
rect 16380 47966 16382 48018
rect 16434 47966 16436 48018
rect 16380 47234 16436 47966
rect 16828 47682 16884 48524
rect 18060 49196 18228 49252
rect 18284 50372 18340 50382
rect 17612 48132 17668 48142
rect 17612 48038 17668 48076
rect 18060 48132 18116 49196
rect 18060 48066 18116 48076
rect 18172 49028 18228 49038
rect 18284 49028 18340 50316
rect 18396 49924 18452 51326
rect 21084 51378 21140 52108
rect 21084 51326 21086 51378
rect 21138 51326 21140 51378
rect 21084 51314 21140 51326
rect 18396 49858 18452 49868
rect 18508 50370 18564 50382
rect 18508 50318 18510 50370
rect 18562 50318 18564 50370
rect 18508 49252 18564 50318
rect 19836 50204 20100 50214
rect 19892 50148 19940 50204
rect 19996 50148 20044 50204
rect 19836 50138 20100 50148
rect 18732 49252 18788 49262
rect 18508 49250 18788 49252
rect 18508 49198 18734 49250
rect 18786 49198 18788 49250
rect 18508 49196 18788 49198
rect 18732 49186 18788 49196
rect 18172 49026 18340 49028
rect 18172 48974 18174 49026
rect 18226 48974 18340 49026
rect 18172 48972 18340 48974
rect 19068 49138 19124 49150
rect 19068 49086 19070 49138
rect 19122 49086 19124 49138
rect 19068 49028 19124 49086
rect 18172 48242 18228 48972
rect 19068 48962 19124 48972
rect 20412 48916 20468 48926
rect 20412 48822 20468 48860
rect 20524 48914 20580 48926
rect 20524 48862 20526 48914
rect 20578 48862 20580 48914
rect 18172 48190 18174 48242
rect 18226 48190 18228 48242
rect 17500 48020 17556 48030
rect 16828 47630 16830 47682
rect 16882 47630 16884 47682
rect 16828 47570 16884 47630
rect 16828 47518 16830 47570
rect 16882 47518 16884 47570
rect 16828 47506 16884 47518
rect 17164 48018 17556 48020
rect 17164 47966 17502 48018
rect 17554 47966 17556 48018
rect 17164 47964 17556 47966
rect 17164 47460 17220 47964
rect 17500 47954 17556 47964
rect 18172 47796 18228 48190
rect 18396 48802 18452 48814
rect 18396 48750 18398 48802
rect 18450 48750 18452 48802
rect 17164 47366 17220 47404
rect 17388 47740 18228 47796
rect 18284 47908 18340 47918
rect 17276 47348 17332 47358
rect 17388 47348 17444 47740
rect 18284 47684 18340 47852
rect 18172 47628 18340 47684
rect 18396 47684 18452 48750
rect 18956 48802 19012 48814
rect 18956 48750 18958 48802
rect 19010 48750 19012 48802
rect 18620 48242 18676 48254
rect 18620 48190 18622 48242
rect 18674 48190 18676 48242
rect 18620 48132 18676 48190
rect 18620 48066 18676 48076
rect 18732 48130 18788 48142
rect 18732 48078 18734 48130
rect 18786 48078 18788 48130
rect 18620 47796 18676 47806
rect 18508 47684 18564 47694
rect 18396 47628 18508 47684
rect 18172 47570 18228 47628
rect 18508 47590 18564 47628
rect 18172 47518 18174 47570
rect 18226 47518 18228 47570
rect 18172 47506 18228 47518
rect 18284 47460 18340 47470
rect 18620 47460 18676 47740
rect 18284 47366 18340 47404
rect 18396 47404 18676 47460
rect 17276 47346 17444 47348
rect 17276 47294 17278 47346
rect 17330 47294 17444 47346
rect 17276 47292 17444 47294
rect 17276 47282 17332 47292
rect 16380 47182 16382 47234
rect 16434 47182 16436 47234
rect 16380 46452 16436 47182
rect 17500 47236 17556 47246
rect 17500 47234 17668 47236
rect 17500 47182 17502 47234
rect 17554 47182 17668 47234
rect 17500 47180 17668 47182
rect 17500 47170 17556 47180
rect 16380 46386 16436 46396
rect 16268 45726 16270 45778
rect 16322 45726 16324 45778
rect 16268 45714 16324 45726
rect 16492 45890 16548 45902
rect 16492 45838 16494 45890
rect 16546 45838 16548 45890
rect 16492 45780 16548 45838
rect 16716 45892 16772 45902
rect 16716 45798 16772 45836
rect 17388 45892 17444 45902
rect 16492 45714 16548 45724
rect 16156 45666 16212 45678
rect 16156 45614 16158 45666
rect 16210 45614 16212 45666
rect 16156 44434 16212 45614
rect 17388 45666 17444 45836
rect 17388 45614 17390 45666
rect 17442 45614 17444 45666
rect 16156 44382 16158 44434
rect 16210 44382 16212 44434
rect 16156 44370 16212 44382
rect 16268 44996 16324 45006
rect 16268 43988 16324 44940
rect 17388 44884 17444 45614
rect 17388 44818 17444 44828
rect 17500 44436 17556 44446
rect 17052 44380 17500 44436
rect 15932 40462 15934 40514
rect 15986 40462 15988 40514
rect 15932 40450 15988 40462
rect 16156 40740 16212 40750
rect 16156 40514 16212 40684
rect 16156 40462 16158 40514
rect 16210 40462 16212 40514
rect 15820 38332 15988 38388
rect 15708 38322 15764 38332
rect 15932 38164 15988 38332
rect 15820 38108 15988 38164
rect 15596 37998 15598 38050
rect 15650 37998 15652 38050
rect 15596 37986 15652 37998
rect 15708 38052 15764 38062
rect 15708 37828 15764 37996
rect 15708 37734 15764 37772
rect 15820 37604 15876 38108
rect 15372 37266 15540 37268
rect 15372 37214 15374 37266
rect 15426 37214 15540 37266
rect 15372 37212 15540 37214
rect 15708 37548 15876 37604
rect 15932 37938 15988 37950
rect 15932 37886 15934 37938
rect 15986 37886 15988 37938
rect 15372 37202 15428 37212
rect 14924 37154 14980 37166
rect 14924 37102 14926 37154
rect 14978 37102 14980 37154
rect 14924 36708 14980 37102
rect 14924 36642 14980 36652
rect 15036 35924 15092 35934
rect 15036 35830 15092 35868
rect 14812 35812 14868 35822
rect 14812 35810 14980 35812
rect 14812 35758 14814 35810
rect 14866 35758 14980 35810
rect 14812 35756 14980 35758
rect 14812 35746 14868 35756
rect 14700 35698 14756 35710
rect 14700 35646 14702 35698
rect 14754 35646 14756 35698
rect 14700 35028 14756 35646
rect 14924 35364 14980 35756
rect 14924 35298 14980 35308
rect 15372 35588 15428 35598
rect 15372 35364 15428 35532
rect 15372 35298 15428 35308
rect 14700 34962 14756 34972
rect 14924 34914 14980 34926
rect 14924 34862 14926 34914
rect 14978 34862 14980 34914
rect 14812 34802 14868 34814
rect 14812 34750 14814 34802
rect 14866 34750 14868 34802
rect 14364 34130 14644 34132
rect 14364 34078 14366 34130
rect 14418 34078 14644 34130
rect 14364 34076 14644 34078
rect 14700 34692 14756 34702
rect 14700 34242 14756 34636
rect 14812 34468 14868 34750
rect 14812 34402 14868 34412
rect 14700 34190 14702 34242
rect 14754 34190 14756 34242
rect 14364 33570 14420 34076
rect 14700 33908 14756 34190
rect 14924 34020 14980 34862
rect 14924 33954 14980 33964
rect 15036 34356 15092 34366
rect 14700 33842 14756 33852
rect 15036 33684 15092 34300
rect 15260 34132 15316 34142
rect 15596 34132 15652 34142
rect 15260 34130 15596 34132
rect 15260 34078 15262 34130
rect 15314 34078 15596 34130
rect 15260 34076 15596 34078
rect 15260 34066 15316 34076
rect 15036 33628 15428 33684
rect 14364 33518 14366 33570
rect 14418 33518 14420 33570
rect 14364 33506 14420 33518
rect 14588 33572 14644 33582
rect 13916 33404 14196 33460
rect 14588 33458 14644 33516
rect 14588 33406 14590 33458
rect 14642 33406 14644 33458
rect 13692 33124 13748 33134
rect 13468 32734 13470 32786
rect 13522 32734 13524 32786
rect 13468 32340 13524 32734
rect 13580 33122 13748 33124
rect 13580 33070 13694 33122
rect 13746 33070 13748 33122
rect 13580 33068 13748 33070
rect 13580 32564 13636 33068
rect 13692 33058 13748 33068
rect 13916 32900 13972 33404
rect 14028 33236 14084 33246
rect 14084 33180 14196 33236
rect 14028 33170 14084 33180
rect 14140 33122 14196 33180
rect 14140 33070 14142 33122
rect 14194 33070 14196 33122
rect 14140 33058 14196 33070
rect 13916 32844 14196 32900
rect 13916 32676 13972 32686
rect 13916 32582 13972 32620
rect 13580 32498 13636 32508
rect 13468 32284 13972 32340
rect 13356 32050 13412 32060
rect 12908 30940 13300 30996
rect 13356 31892 13412 31902
rect 13356 30994 13412 31836
rect 13468 31778 13524 31790
rect 13468 31726 13470 31778
rect 13522 31726 13524 31778
rect 13468 31108 13524 31726
rect 13916 31780 13972 32284
rect 13468 31042 13524 31052
rect 13804 31332 13860 31342
rect 13356 30942 13358 30994
rect 13410 30942 13412 30994
rect 12684 30716 12852 30772
rect 12572 30046 12574 30098
rect 12626 30046 12628 30098
rect 12460 29428 12516 29438
rect 12236 29426 12516 29428
rect 12236 29374 12462 29426
rect 12514 29374 12516 29426
rect 12236 29372 12516 29374
rect 12124 29314 12180 29372
rect 12124 29262 12126 29314
rect 12178 29262 12180 29314
rect 12124 29250 12180 29262
rect 11900 28702 11902 28754
rect 11954 28702 11956 28754
rect 11900 28690 11956 28702
rect 12236 28868 12292 28878
rect 12236 28754 12292 28812
rect 12236 28702 12238 28754
rect 12290 28702 12292 28754
rect 12236 28690 12292 28702
rect 11340 28590 11342 28642
rect 11394 28590 11396 28642
rect 11340 28578 11396 28590
rect 11564 28084 11620 28094
rect 11564 27990 11620 28028
rect 12236 28084 12292 28094
rect 12124 27860 12180 27870
rect 12124 27766 12180 27804
rect 12236 27300 12292 28028
rect 12124 27244 12292 27300
rect 12348 27970 12404 27982
rect 12348 27918 12350 27970
rect 12402 27918 12404 27970
rect 12348 27300 12404 27918
rect 12124 26908 12180 27244
rect 12236 27076 12292 27114
rect 12236 27010 12292 27020
rect 11788 26852 11844 26862
rect 12124 26852 12292 26908
rect 11452 26628 11508 26638
rect 11340 26292 11396 26302
rect 11228 26290 11396 26292
rect 11228 26238 11342 26290
rect 11394 26238 11396 26290
rect 11228 26236 11396 26238
rect 11340 26226 11396 26236
rect 11452 26068 11508 26572
rect 11004 25890 11060 25900
rect 11228 26012 11508 26068
rect 10444 25506 10500 25518
rect 10444 25454 10446 25506
rect 10498 25454 10500 25506
rect 10444 25396 10500 25454
rect 11004 25508 11060 25518
rect 11004 25414 11060 25452
rect 10444 25330 10500 25340
rect 10780 25396 10836 25406
rect 10780 25302 10836 25340
rect 11228 24946 11284 26012
rect 11788 25506 11844 26796
rect 12012 26628 12068 26638
rect 11900 26292 11956 26302
rect 11900 26198 11956 26236
rect 11788 25454 11790 25506
rect 11842 25454 11844 25506
rect 11788 25442 11844 25454
rect 11900 25508 11956 25518
rect 11900 25414 11956 25452
rect 12012 25506 12068 26572
rect 12236 26290 12292 26852
rect 12236 26238 12238 26290
rect 12290 26238 12292 26290
rect 12236 26226 12292 26238
rect 12012 25454 12014 25506
rect 12066 25454 12068 25506
rect 12012 25442 12068 25454
rect 12348 25506 12404 27244
rect 12348 25454 12350 25506
rect 12402 25454 12404 25506
rect 11228 24894 11230 24946
rect 11282 24894 11284 24946
rect 11228 24882 11284 24894
rect 11340 25282 11396 25294
rect 11340 25230 11342 25282
rect 11394 25230 11396 25282
rect 11340 24164 11396 25230
rect 11676 24948 11732 24986
rect 11676 24882 11732 24892
rect 12348 24948 12404 25454
rect 12460 25284 12516 29372
rect 12572 28532 12628 30046
rect 12684 29988 12740 29998
rect 12684 29316 12740 29932
rect 12684 29250 12740 29260
rect 12684 28756 12740 28766
rect 12684 28662 12740 28700
rect 12572 28466 12628 28476
rect 12684 27860 12740 27870
rect 12684 27186 12740 27804
rect 12684 27134 12686 27186
rect 12738 27134 12740 27186
rect 12684 27122 12740 27134
rect 12796 26908 12852 30716
rect 12908 30210 12964 30940
rect 13356 30930 13412 30942
rect 12908 30158 12910 30210
rect 12962 30158 12964 30210
rect 12908 30146 12964 30158
rect 13020 30772 13076 30782
rect 13020 28082 13076 30716
rect 13692 30100 13748 30110
rect 13580 29986 13636 29998
rect 13580 29934 13582 29986
rect 13634 29934 13636 29986
rect 13580 29876 13636 29934
rect 13356 29764 13412 29774
rect 13356 29426 13412 29708
rect 13356 29374 13358 29426
rect 13410 29374 13412 29426
rect 13132 29204 13188 29214
rect 13132 29202 13300 29204
rect 13132 29150 13134 29202
rect 13186 29150 13300 29202
rect 13132 29148 13300 29150
rect 13132 29138 13188 29148
rect 13020 28030 13022 28082
rect 13074 28030 13076 28082
rect 13020 28018 13076 28030
rect 13244 28532 13300 29148
rect 13356 28756 13412 29374
rect 13356 28690 13412 28700
rect 13580 28644 13636 29820
rect 13692 29538 13748 30044
rect 13692 29486 13694 29538
rect 13746 29486 13748 29538
rect 13692 29316 13748 29486
rect 13804 29540 13860 31276
rect 13916 31106 13972 31724
rect 14028 32004 14084 32014
rect 14028 31778 14084 31948
rect 14028 31726 14030 31778
rect 14082 31726 14084 31778
rect 14028 31714 14084 31726
rect 13916 31054 13918 31106
rect 13970 31054 13972 31106
rect 13916 31042 13972 31054
rect 14140 31218 14196 32844
rect 14252 32676 14308 32686
rect 14252 32582 14308 32620
rect 14588 32676 14644 33406
rect 14588 32610 14644 32620
rect 14924 33570 14980 33582
rect 14924 33518 14926 33570
rect 14978 33518 14980 33570
rect 14924 33124 14980 33518
rect 15036 33124 15092 33134
rect 14924 33068 15036 33124
rect 14700 32450 14756 32462
rect 14700 32398 14702 32450
rect 14754 32398 14756 32450
rect 14588 31666 14644 31678
rect 14588 31614 14590 31666
rect 14642 31614 14644 31666
rect 14588 31332 14644 31614
rect 14140 31166 14142 31218
rect 14194 31166 14196 31218
rect 14140 30996 14196 31166
rect 14252 31276 14644 31332
rect 14252 31108 14308 31276
rect 14476 31108 14532 31118
rect 14252 31042 14308 31052
rect 14364 31052 14476 31108
rect 14140 30930 14196 30940
rect 14364 30994 14420 31052
rect 14476 31042 14532 31052
rect 14364 30942 14366 30994
rect 14418 30942 14420 30994
rect 14252 30882 14308 30894
rect 14252 30830 14254 30882
rect 14306 30830 14308 30882
rect 14140 30660 14196 30670
rect 14140 29988 14196 30604
rect 14252 30212 14308 30830
rect 14364 30434 14420 30942
rect 14364 30382 14366 30434
rect 14418 30382 14420 30434
rect 14364 30370 14420 30382
rect 14588 30996 14644 31006
rect 14700 30996 14756 32398
rect 14812 31780 14868 31790
rect 14812 31686 14868 31724
rect 14588 30994 14756 30996
rect 14588 30942 14590 30994
rect 14642 30942 14756 30994
rect 14588 30940 14756 30942
rect 14588 30436 14644 30940
rect 14588 30370 14644 30380
rect 14700 30434 14756 30446
rect 14700 30382 14702 30434
rect 14754 30382 14756 30434
rect 14700 30324 14756 30382
rect 14700 30322 14868 30324
rect 14700 30270 14702 30322
rect 14754 30270 14868 30322
rect 14700 30268 14868 30270
rect 14700 30258 14756 30268
rect 14252 30156 14644 30212
rect 14252 29988 14308 29998
rect 14140 29986 14308 29988
rect 14140 29934 14254 29986
rect 14306 29934 14308 29986
rect 14140 29932 14308 29934
rect 14252 29922 14308 29932
rect 14588 29764 14644 30156
rect 14588 29708 14756 29764
rect 13916 29540 13972 29550
rect 13804 29538 13972 29540
rect 13804 29486 13918 29538
rect 13970 29486 13972 29538
rect 13804 29484 13972 29486
rect 13916 29474 13972 29484
rect 14700 29538 14756 29708
rect 14700 29486 14702 29538
rect 14754 29486 14756 29538
rect 14700 29474 14756 29486
rect 14364 29426 14420 29438
rect 14364 29374 14366 29426
rect 14418 29374 14420 29426
rect 14364 29316 14420 29374
rect 13692 29250 13748 29260
rect 13916 29260 14420 29316
rect 14588 29426 14644 29438
rect 14588 29374 14590 29426
rect 14642 29374 14644 29426
rect 13804 29204 13860 29214
rect 13916 29204 13972 29260
rect 13804 29202 13972 29204
rect 13804 29150 13806 29202
rect 13858 29150 13972 29202
rect 13804 29148 13972 29150
rect 13804 29138 13860 29148
rect 14588 28980 14644 29374
rect 14812 29428 14868 30268
rect 14924 30100 14980 33068
rect 15036 33030 15092 33068
rect 15036 32900 15092 32910
rect 15036 31778 15092 32844
rect 15260 32450 15316 32462
rect 15260 32398 15262 32450
rect 15314 32398 15316 32450
rect 15260 32004 15316 32398
rect 15260 31938 15316 31948
rect 15036 31726 15038 31778
rect 15090 31726 15092 31778
rect 15036 30660 15092 31726
rect 15148 31890 15204 31902
rect 15148 31838 15150 31890
rect 15202 31838 15204 31890
rect 15148 31780 15204 31838
rect 15148 31724 15316 31780
rect 15260 31668 15316 31724
rect 15260 31602 15316 31612
rect 15148 31554 15204 31566
rect 15148 31502 15150 31554
rect 15202 31502 15204 31554
rect 15148 31444 15204 31502
rect 15372 31444 15428 33628
rect 15484 33460 15540 33470
rect 15484 33366 15540 33404
rect 15148 31388 15428 31444
rect 15148 31220 15204 31230
rect 15372 31220 15428 31230
rect 15148 31218 15372 31220
rect 15148 31166 15150 31218
rect 15202 31166 15372 31218
rect 15148 31164 15372 31166
rect 15148 31154 15204 31164
rect 15372 31154 15428 31164
rect 15484 31108 15540 31118
rect 15484 31014 15540 31052
rect 15036 30594 15092 30604
rect 15260 30996 15316 31006
rect 15260 30322 15316 30940
rect 15260 30270 15262 30322
rect 15314 30270 15316 30322
rect 15260 30258 15316 30270
rect 14924 30034 14980 30044
rect 15148 29988 15204 29998
rect 15148 29650 15204 29932
rect 15148 29598 15150 29650
rect 15202 29598 15204 29650
rect 15148 29586 15204 29598
rect 14812 29362 14868 29372
rect 15596 29314 15652 34076
rect 15708 31780 15764 37548
rect 15932 37492 15988 37886
rect 16156 37604 16212 40462
rect 16268 39396 16324 43932
rect 16380 44322 16436 44334
rect 16380 44270 16382 44322
rect 16434 44270 16436 44322
rect 16380 43764 16436 44270
rect 16604 44324 16660 44334
rect 16604 44230 16660 44268
rect 16828 44324 16884 44334
rect 16828 44230 16884 44268
rect 16380 43698 16436 43708
rect 16604 43540 16660 43550
rect 16492 43484 16604 43540
rect 16380 41188 16436 41198
rect 16380 40626 16436 41132
rect 16380 40574 16382 40626
rect 16434 40574 16436 40626
rect 16380 40562 16436 40574
rect 16380 39844 16436 39854
rect 16380 39618 16436 39788
rect 16380 39566 16382 39618
rect 16434 39566 16436 39618
rect 16380 39554 16436 39566
rect 16268 39340 16436 39396
rect 16268 38722 16324 38734
rect 16268 38670 16270 38722
rect 16322 38670 16324 38722
rect 16268 38052 16324 38670
rect 16380 38276 16436 39340
rect 16492 39284 16548 43484
rect 16604 43474 16660 43484
rect 16716 42756 16772 42766
rect 16716 42194 16772 42700
rect 17052 42756 17108 44380
rect 17500 44322 17556 44380
rect 17500 44270 17502 44322
rect 17554 44270 17556 44322
rect 17500 44258 17556 44270
rect 17388 44212 17444 44222
rect 17388 44118 17444 44156
rect 17276 44100 17332 44110
rect 17276 44006 17332 44044
rect 17612 43988 17668 47180
rect 18172 47234 18228 47246
rect 18172 47182 18174 47234
rect 18226 47182 18228 47234
rect 18172 47124 18228 47182
rect 18172 47058 18228 47068
rect 17836 45780 17892 45790
rect 17836 45686 17892 45724
rect 17724 45108 17780 45118
rect 17724 44100 17780 45052
rect 17724 44034 17780 44044
rect 17388 43932 17668 43988
rect 17388 43650 17444 43932
rect 17500 43764 17556 43774
rect 17500 43670 17556 43708
rect 17388 43598 17390 43650
rect 17442 43598 17444 43650
rect 17388 43586 17444 43598
rect 17612 43652 17668 43662
rect 17612 43558 17668 43596
rect 17836 43540 17892 43550
rect 17724 43538 17892 43540
rect 17724 43486 17838 43538
rect 17890 43486 17892 43538
rect 17724 43484 17892 43486
rect 17052 42690 17108 42700
rect 17612 42756 17668 42766
rect 17612 42662 17668 42700
rect 16716 42142 16718 42194
rect 16770 42142 16772 42194
rect 16716 42130 16772 42142
rect 16604 41972 16660 41982
rect 16604 41878 16660 41916
rect 16716 41746 16772 41758
rect 16716 41694 16718 41746
rect 16770 41694 16772 41746
rect 16604 40402 16660 40414
rect 16604 40350 16606 40402
rect 16658 40350 16660 40402
rect 16604 40068 16660 40350
rect 16604 40002 16660 40012
rect 16716 39844 16772 41694
rect 17724 41412 17780 43484
rect 17836 43474 17892 43484
rect 18172 43540 18228 43550
rect 18172 43538 18340 43540
rect 18172 43486 18174 43538
rect 18226 43486 18340 43538
rect 18172 43484 18340 43486
rect 18172 43474 18228 43484
rect 18060 42754 18116 42766
rect 18060 42702 18062 42754
rect 18114 42702 18116 42754
rect 18060 42532 18116 42702
rect 17836 42420 17892 42430
rect 17836 42082 17892 42364
rect 17836 42030 17838 42082
rect 17890 42030 17892 42082
rect 17836 42018 17892 42030
rect 17948 42082 18004 42094
rect 17948 42030 17950 42082
rect 18002 42030 18004 42082
rect 16604 39788 16772 39844
rect 16940 41356 17780 41412
rect 17948 41972 18004 42030
rect 18060 42084 18116 42476
rect 18060 42018 18116 42028
rect 16604 39396 16660 39788
rect 16604 39340 16772 39396
rect 16492 39228 16660 39284
rect 16380 38210 16436 38220
rect 16492 38388 16548 38398
rect 16492 38052 16548 38332
rect 16604 38274 16660 39228
rect 16604 38222 16606 38274
rect 16658 38222 16660 38274
rect 16604 38210 16660 38222
rect 16492 37996 16660 38052
rect 16268 37986 16324 37996
rect 16380 37828 16436 37838
rect 16380 37734 16436 37772
rect 16492 37604 16548 37614
rect 16156 37548 16436 37604
rect 15820 37436 15988 37492
rect 15820 37378 15876 37436
rect 15820 37326 15822 37378
rect 15874 37326 15876 37378
rect 15820 37314 15876 37326
rect 16156 37380 16212 37390
rect 16044 37266 16100 37278
rect 16044 37214 16046 37266
rect 16098 37214 16100 37266
rect 16044 35924 16100 37214
rect 16156 37154 16212 37324
rect 16268 37268 16324 37278
rect 16268 37174 16324 37212
rect 16156 37102 16158 37154
rect 16210 37102 16212 37154
rect 16156 37090 16212 37102
rect 16380 36260 16436 37548
rect 16492 37380 16548 37548
rect 16492 37286 16548 37324
rect 16604 37044 16660 37996
rect 16380 36194 16436 36204
rect 16492 36988 16660 37044
rect 16044 35858 16100 35868
rect 16268 35588 16324 35598
rect 15932 35028 15988 35038
rect 15820 34802 15876 34814
rect 15820 34750 15822 34802
rect 15874 34750 15876 34802
rect 15820 34354 15876 34750
rect 15820 34302 15822 34354
rect 15874 34302 15876 34354
rect 15820 34290 15876 34302
rect 15932 34242 15988 34972
rect 15932 34190 15934 34242
rect 15986 34190 15988 34242
rect 15932 33236 15988 34190
rect 15932 33170 15988 33180
rect 16044 34914 16100 34926
rect 16044 34862 16046 34914
rect 16098 34862 16100 34914
rect 16044 31892 16100 34862
rect 16156 34130 16212 34142
rect 16156 34078 16158 34130
rect 16210 34078 16212 34130
rect 16156 33570 16212 34078
rect 16156 33518 16158 33570
rect 16210 33518 16212 33570
rect 16156 33506 16212 33518
rect 15932 31836 16100 31892
rect 16156 33236 16212 33246
rect 16156 32004 16212 33180
rect 16268 32900 16324 35532
rect 16380 33572 16436 33582
rect 16492 33572 16548 36988
rect 16716 34804 16772 39340
rect 16940 38836 16996 41356
rect 16940 35812 16996 38780
rect 17164 41186 17220 41198
rect 17164 41134 17166 41186
rect 17218 41134 17220 41186
rect 17164 38668 17220 41134
rect 17612 41188 17668 41198
rect 17612 41094 17668 41132
rect 17500 40740 17556 40750
rect 17500 40516 17556 40684
rect 17500 40402 17556 40460
rect 17500 40350 17502 40402
rect 17554 40350 17556 40402
rect 17500 40338 17556 40350
rect 17724 40514 17780 40526
rect 17724 40462 17726 40514
rect 17778 40462 17780 40514
rect 17724 40180 17780 40462
rect 17724 40114 17780 40124
rect 17388 39732 17444 39742
rect 17388 39618 17444 39676
rect 17388 39566 17390 39618
rect 17442 39566 17444 39618
rect 17388 39554 17444 39566
rect 17052 38612 17220 38668
rect 17052 36708 17108 38612
rect 17164 38052 17220 38062
rect 17836 38052 17892 38062
rect 17164 38050 17444 38052
rect 17164 37998 17166 38050
rect 17218 37998 17444 38050
rect 17164 37996 17444 37998
rect 17164 37986 17220 37996
rect 17276 37826 17332 37838
rect 17276 37774 17278 37826
rect 17330 37774 17332 37826
rect 17276 37492 17332 37774
rect 17276 37426 17332 37436
rect 17388 37268 17444 37996
rect 17836 37958 17892 37996
rect 17724 37940 17780 37950
rect 17724 37846 17780 37884
rect 17500 37828 17556 37838
rect 17500 37826 17668 37828
rect 17500 37774 17502 37826
rect 17554 37774 17668 37826
rect 17500 37772 17668 37774
rect 17500 37762 17556 37772
rect 17052 36652 17332 36708
rect 16940 35756 17220 35812
rect 16940 34916 16996 34926
rect 16940 34822 16996 34860
rect 16604 34748 16772 34804
rect 16828 34804 16884 34814
rect 16604 33684 16660 34748
rect 16828 34710 16884 34748
rect 17052 34244 17108 34254
rect 16716 34132 16772 34142
rect 16716 34038 16772 34076
rect 16604 33618 16660 33628
rect 16940 33796 16996 33806
rect 16380 33570 16548 33572
rect 16380 33518 16382 33570
rect 16434 33518 16548 33570
rect 16380 33516 16548 33518
rect 16380 33122 16436 33516
rect 16380 33070 16382 33122
rect 16434 33070 16436 33122
rect 16380 33012 16436 33070
rect 16940 33124 16996 33740
rect 17052 33684 17108 34188
rect 17052 33618 17108 33628
rect 17164 33458 17220 35756
rect 17276 35026 17332 36652
rect 17276 34974 17278 35026
rect 17330 34974 17332 35026
rect 17276 34962 17332 34974
rect 17388 33908 17444 37212
rect 17500 37604 17556 37614
rect 17500 37266 17556 37548
rect 17500 37214 17502 37266
rect 17554 37214 17556 37266
rect 17500 36372 17556 37214
rect 17500 36278 17556 36316
rect 17612 36036 17668 37772
rect 17836 37380 17892 37390
rect 17948 37380 18004 41916
rect 18172 41972 18228 41982
rect 18172 41878 18228 41916
rect 18284 40740 18340 43484
rect 18396 41298 18452 47404
rect 18620 47124 18676 47134
rect 18620 45220 18676 47068
rect 18508 45164 18676 45220
rect 18508 41972 18564 45164
rect 18620 44994 18676 45006
rect 18620 44942 18622 44994
rect 18674 44942 18676 44994
rect 18620 44548 18676 44942
rect 18620 44482 18676 44492
rect 18732 44212 18788 48078
rect 18956 47908 19012 48750
rect 19628 48802 19684 48814
rect 19628 48750 19630 48802
rect 19682 48750 19684 48802
rect 19292 48354 19348 48366
rect 19292 48302 19294 48354
rect 19346 48302 19348 48354
rect 19180 48132 19236 48142
rect 19012 47852 19124 47908
rect 18956 47842 19012 47852
rect 18956 47684 19012 47694
rect 18956 47346 19012 47628
rect 18956 47294 18958 47346
rect 19010 47294 19012 47346
rect 18956 47282 19012 47294
rect 18732 44146 18788 44156
rect 19068 45330 19124 47852
rect 19180 47458 19236 48076
rect 19292 47682 19348 48302
rect 19628 48356 19684 48750
rect 20188 48802 20244 48814
rect 20188 48750 20190 48802
rect 20242 48750 20244 48802
rect 19836 48636 20100 48646
rect 19892 48580 19940 48636
rect 19996 48580 20044 48636
rect 19836 48570 20100 48580
rect 20188 48468 20244 48750
rect 19628 48262 19684 48300
rect 20076 48412 20244 48468
rect 20076 48242 20132 48412
rect 20076 48190 20078 48242
rect 20130 48190 20132 48242
rect 20076 48178 20132 48190
rect 20524 48244 20580 48862
rect 20524 48178 20580 48188
rect 20300 48130 20356 48142
rect 20300 48078 20302 48130
rect 20354 48078 20356 48130
rect 19292 47630 19294 47682
rect 19346 47630 19348 47682
rect 19292 47618 19348 47630
rect 20076 47684 20132 47694
rect 20132 47628 20244 47684
rect 20076 47618 20132 47628
rect 19180 47406 19182 47458
rect 19234 47406 19236 47458
rect 19180 47394 19236 47406
rect 19516 47460 19572 47470
rect 19740 47460 19796 47470
rect 19516 47458 19796 47460
rect 19516 47406 19518 47458
rect 19570 47406 19742 47458
rect 19794 47406 19796 47458
rect 19516 47404 19796 47406
rect 19516 47394 19572 47404
rect 19628 46564 19684 47404
rect 19740 47394 19796 47404
rect 20076 47460 20132 47470
rect 20076 47236 20132 47404
rect 20188 47348 20244 47628
rect 20300 47460 20356 48078
rect 20300 47404 20580 47460
rect 20188 47292 20356 47348
rect 20076 47180 20244 47236
rect 19836 47068 20100 47078
rect 19892 47012 19940 47068
rect 19996 47012 20044 47068
rect 19836 47002 20100 47012
rect 20188 46900 20244 47180
rect 19964 46844 20244 46900
rect 20300 47234 20356 47292
rect 20300 47182 20302 47234
rect 20354 47182 20356 47234
rect 19964 46786 20020 46844
rect 19964 46734 19966 46786
rect 20018 46734 20020 46786
rect 19964 46722 20020 46734
rect 19628 46498 19684 46508
rect 20076 46676 20132 46686
rect 19964 45892 20020 45902
rect 19068 45278 19070 45330
rect 19122 45278 19124 45330
rect 18732 43650 18788 43662
rect 18732 43598 18734 43650
rect 18786 43598 18788 43650
rect 18620 43540 18676 43550
rect 18620 43446 18676 43484
rect 18732 42980 18788 43598
rect 19068 43652 19124 45278
rect 19180 45890 20020 45892
rect 19180 45838 19966 45890
rect 20018 45838 20020 45890
rect 19180 45836 20020 45838
rect 19180 44210 19236 45836
rect 19404 45218 19460 45836
rect 19964 45826 20020 45836
rect 20076 45890 20132 46620
rect 20300 46674 20356 47182
rect 20300 46622 20302 46674
rect 20354 46622 20356 46674
rect 20300 46610 20356 46622
rect 20412 47234 20468 47246
rect 20412 47182 20414 47234
rect 20466 47182 20468 47234
rect 20076 45838 20078 45890
rect 20130 45838 20132 45890
rect 20076 45826 20132 45838
rect 20300 46450 20356 46462
rect 20300 46398 20302 46450
rect 20354 46398 20356 46450
rect 20300 45892 20356 46398
rect 20300 45826 20356 45836
rect 19740 45668 19796 45678
rect 19628 45666 19796 45668
rect 19628 45614 19742 45666
rect 19794 45614 19796 45666
rect 19628 45612 19796 45614
rect 19628 45556 19684 45612
rect 19740 45602 19796 45612
rect 20188 45556 20244 45566
rect 19628 45490 19684 45500
rect 19836 45500 20100 45510
rect 19892 45444 19940 45500
rect 19996 45444 20044 45500
rect 19836 45434 20100 45444
rect 19404 45166 19406 45218
rect 19458 45166 19460 45218
rect 19404 45154 19460 45166
rect 19628 45218 19684 45230
rect 19628 45166 19630 45218
rect 19682 45166 19684 45218
rect 19628 44436 19684 45166
rect 19964 45106 20020 45118
rect 19964 45054 19966 45106
rect 20018 45054 20020 45106
rect 19964 44660 20020 45054
rect 20188 44772 20244 45500
rect 20300 44996 20356 45006
rect 20300 44902 20356 44940
rect 20188 44716 20356 44772
rect 19964 44594 20020 44604
rect 19628 44370 19684 44380
rect 19180 44158 19182 44210
rect 19234 44158 19236 44210
rect 19180 44146 19236 44158
rect 19852 44212 19908 44222
rect 19852 44118 19908 44156
rect 19068 43586 19124 43596
rect 19292 44100 19348 44110
rect 18732 42914 18788 42924
rect 18732 42644 18788 42654
rect 18620 41972 18676 41982
rect 18508 41970 18676 41972
rect 18508 41918 18622 41970
rect 18674 41918 18676 41970
rect 18508 41916 18676 41918
rect 18620 41906 18676 41916
rect 18508 41748 18564 41758
rect 18508 41746 18676 41748
rect 18508 41694 18510 41746
rect 18562 41694 18676 41746
rect 18508 41692 18676 41694
rect 18508 41682 18564 41692
rect 18396 41246 18398 41298
rect 18450 41246 18452 41298
rect 18396 41234 18452 41246
rect 18284 40674 18340 40684
rect 18172 40628 18228 40638
rect 18172 40534 18228 40572
rect 18508 40292 18564 40302
rect 18508 40198 18564 40236
rect 18172 39508 18228 39518
rect 18172 38948 18228 39452
rect 18620 39396 18676 41692
rect 18732 41074 18788 42588
rect 18844 41748 18900 41758
rect 18844 41654 18900 41692
rect 18956 41748 19012 41758
rect 18956 41746 19124 41748
rect 18956 41694 18958 41746
rect 19010 41694 19124 41746
rect 18956 41692 19124 41694
rect 18956 41682 19012 41692
rect 18732 41022 18734 41074
rect 18786 41022 18788 41074
rect 18732 41010 18788 41022
rect 18732 40628 18788 40638
rect 18732 40514 18788 40572
rect 18732 40462 18734 40514
rect 18786 40462 18788 40514
rect 18732 40450 18788 40462
rect 18844 40402 18900 40414
rect 18844 40350 18846 40402
rect 18898 40350 18900 40402
rect 18620 39340 18788 39396
rect 18172 38882 18228 38892
rect 18060 38722 18116 38734
rect 18060 38670 18062 38722
rect 18114 38670 18116 38722
rect 18060 38668 18116 38670
rect 18620 38722 18676 38734
rect 18620 38670 18622 38722
rect 18674 38670 18676 38722
rect 18620 38668 18676 38670
rect 18060 38612 18676 38668
rect 18284 38050 18340 38062
rect 18284 37998 18286 38050
rect 18338 37998 18340 38050
rect 18284 37604 18340 37998
rect 18284 37538 18340 37548
rect 18396 37492 18452 38612
rect 18732 38276 18788 39340
rect 18620 38220 18788 38276
rect 18844 38276 18900 40350
rect 19068 40402 19124 41692
rect 19068 40350 19070 40402
rect 19122 40350 19124 40402
rect 19068 40338 19124 40350
rect 18956 39618 19012 39630
rect 18956 39566 18958 39618
rect 19010 39566 19012 39618
rect 18956 39284 19012 39566
rect 18956 39218 19012 39228
rect 19068 38722 19124 38734
rect 19068 38670 19070 38722
rect 19122 38670 19124 38722
rect 19068 38500 19124 38670
rect 19068 38444 19236 38500
rect 19068 38276 19124 38286
rect 18844 38274 19124 38276
rect 18844 38222 19070 38274
rect 19122 38222 19124 38274
rect 18844 38220 19124 38222
rect 18508 38052 18564 38062
rect 18508 37958 18564 37996
rect 18620 37716 18676 38220
rect 19068 38210 19124 38220
rect 17836 37378 18004 37380
rect 17836 37326 17838 37378
rect 17890 37326 18004 37378
rect 17836 37324 18004 37326
rect 18284 37380 18340 37390
rect 17836 37268 17892 37324
rect 18284 37286 18340 37324
rect 18396 37378 18452 37436
rect 18396 37326 18398 37378
rect 18450 37326 18452 37378
rect 17836 37202 17892 37212
rect 18396 36820 18452 37326
rect 18396 36754 18452 36764
rect 18508 37660 18676 37716
rect 18732 38050 18788 38062
rect 18732 37998 18734 38050
rect 18786 37998 18788 38050
rect 18060 36708 18116 36718
rect 18060 36594 18116 36652
rect 18508 36708 18564 37660
rect 18620 37492 18676 37502
rect 18732 37492 18788 37998
rect 18956 38050 19012 38062
rect 18956 37998 18958 38050
rect 19010 37998 19012 38050
rect 18956 37828 19012 37998
rect 18956 37762 19012 37772
rect 19068 37940 19124 37950
rect 18620 37490 18788 37492
rect 18620 37438 18622 37490
rect 18674 37438 18788 37490
rect 18620 37436 18788 37438
rect 18620 37426 18676 37436
rect 19068 37266 19124 37884
rect 19180 37716 19236 38444
rect 19180 37650 19236 37660
rect 19180 37492 19236 37502
rect 19180 37398 19236 37436
rect 19068 37214 19070 37266
rect 19122 37214 19124 37266
rect 18508 36642 18564 36652
rect 18620 37156 18676 37166
rect 18060 36542 18062 36594
rect 18114 36542 18116 36594
rect 18060 36530 18116 36542
rect 17948 36484 18004 36494
rect 18620 36484 18676 37100
rect 19068 36932 19124 37214
rect 17948 36372 18004 36428
rect 18508 36428 18676 36484
rect 18844 36876 19124 36932
rect 18060 36372 18116 36382
rect 17948 36370 18116 36372
rect 17948 36318 18062 36370
rect 18114 36318 18116 36370
rect 17948 36316 18116 36318
rect 18060 36306 18116 36316
rect 18284 36370 18340 36382
rect 18284 36318 18286 36370
rect 18338 36318 18340 36370
rect 17836 36260 17892 36270
rect 17836 36166 17892 36204
rect 18172 36148 18228 36158
rect 17612 35980 18004 36036
rect 17724 35812 17780 35822
rect 17724 35718 17780 35756
rect 17612 35698 17668 35710
rect 17612 35646 17614 35698
rect 17666 35646 17668 35698
rect 17612 34356 17668 35646
rect 17948 34468 18004 35980
rect 17948 34402 18004 34412
rect 17612 34290 17668 34300
rect 17500 34244 17556 34254
rect 18060 34244 18116 34254
rect 17500 34150 17556 34188
rect 17948 34242 18116 34244
rect 17948 34190 18062 34242
rect 18114 34190 18116 34242
rect 17948 34188 18116 34190
rect 17612 34130 17668 34142
rect 17612 34078 17614 34130
rect 17666 34078 17668 34130
rect 17612 34020 17668 34078
rect 17500 33908 17556 33918
rect 17388 33906 17556 33908
rect 17388 33854 17502 33906
rect 17554 33854 17556 33906
rect 17388 33852 17556 33854
rect 17500 33842 17556 33852
rect 17164 33406 17166 33458
rect 17218 33406 17220 33458
rect 17164 33394 17220 33406
rect 17388 33572 17444 33582
rect 16940 33058 16996 33068
rect 17164 33234 17220 33246
rect 17164 33182 17166 33234
rect 17218 33182 17220 33234
rect 17164 33124 17220 33182
rect 16380 32956 16660 33012
rect 16268 32844 16436 32900
rect 15820 31780 15876 31790
rect 15708 31778 15876 31780
rect 15708 31726 15822 31778
rect 15874 31726 15876 31778
rect 15708 31724 15876 31726
rect 15708 31108 15764 31724
rect 15820 31714 15876 31724
rect 15708 31042 15764 31052
rect 15596 29262 15598 29314
rect 15650 29262 15652 29314
rect 14588 28924 15092 28980
rect 14364 28756 14420 28766
rect 14420 28700 14532 28756
rect 14364 28690 14420 28700
rect 13580 28588 13972 28644
rect 13244 27860 13300 28476
rect 13692 27860 13748 27870
rect 13300 27858 13748 27860
rect 13300 27806 13694 27858
rect 13746 27806 13748 27858
rect 13300 27804 13748 27806
rect 13244 27766 13300 27804
rect 13692 27794 13748 27804
rect 13580 27076 13636 27086
rect 13580 26982 13636 27020
rect 12796 26852 12964 26908
rect 12684 26796 12964 26852
rect 12572 25396 12628 25406
rect 12572 25302 12628 25340
rect 12460 25218 12516 25228
rect 12348 24882 12404 24892
rect 11340 24098 11396 24108
rect 11676 24724 11732 24734
rect 11676 24050 11732 24668
rect 11676 23998 11678 24050
rect 11730 23998 11732 24050
rect 11676 23986 11732 23998
rect 10332 23314 10388 23324
rect 12684 21700 12740 26796
rect 13692 26628 13748 26638
rect 12796 26516 12852 26526
rect 12796 25508 12852 26460
rect 13244 26516 13300 26526
rect 13244 26422 13300 26460
rect 13692 26514 13748 26572
rect 13692 26462 13694 26514
rect 13746 26462 13748 26514
rect 13692 26450 13748 26462
rect 13916 26404 13972 28588
rect 14476 28642 14532 28700
rect 15036 28754 15092 28924
rect 15036 28702 15038 28754
rect 15090 28702 15092 28754
rect 15036 28690 15092 28702
rect 15260 28756 15316 28766
rect 14476 28590 14478 28642
rect 14530 28590 14532 28642
rect 14476 28578 14532 28590
rect 15260 28642 15316 28700
rect 15260 28590 15262 28642
rect 15314 28590 15316 28642
rect 15260 28578 15316 28590
rect 14700 28532 14756 28542
rect 14140 28084 14196 28094
rect 14140 27186 14196 28028
rect 14140 27134 14142 27186
rect 14194 27134 14196 27186
rect 14140 27122 14196 27134
rect 14252 27858 14308 27870
rect 14252 27806 14254 27858
rect 14306 27806 14308 27858
rect 14252 27748 14308 27806
rect 13580 26292 13636 26302
rect 12908 25508 12964 25518
rect 12796 25506 13076 25508
rect 12796 25454 12910 25506
rect 12962 25454 13076 25506
rect 12796 25452 13076 25454
rect 12908 25442 12964 25452
rect 12796 25284 12852 25294
rect 12796 25282 12964 25284
rect 12796 25230 12798 25282
rect 12850 25230 12964 25282
rect 12796 25228 12964 25230
rect 12796 25218 12852 25228
rect 12908 24722 12964 25228
rect 12908 24670 12910 24722
rect 12962 24670 12964 24722
rect 12908 24276 12964 24670
rect 12908 24210 12964 24220
rect 13020 24050 13076 25452
rect 13468 25284 13524 25294
rect 13468 25190 13524 25228
rect 13356 24836 13412 24846
rect 13356 24722 13412 24780
rect 13356 24670 13358 24722
rect 13410 24670 13412 24722
rect 13356 24658 13412 24670
rect 13580 24722 13636 26236
rect 13916 25618 13972 26348
rect 14140 26178 14196 26190
rect 14140 26126 14142 26178
rect 14194 26126 14196 26178
rect 14140 25844 14196 26126
rect 14140 25778 14196 25788
rect 13916 25566 13918 25618
rect 13970 25566 13972 25618
rect 13916 25554 13972 25566
rect 13580 24670 13582 24722
rect 13634 24670 13636 24722
rect 13580 24658 13636 24670
rect 13916 25284 13972 25294
rect 13916 24722 13972 25228
rect 13916 24670 13918 24722
rect 13970 24670 13972 24722
rect 13916 24658 13972 24670
rect 14028 25172 14084 25182
rect 13020 23998 13022 24050
rect 13074 23998 13076 24050
rect 13020 23986 13076 23998
rect 14028 24050 14084 25116
rect 14252 24836 14308 27692
rect 14476 27300 14532 27310
rect 14476 27186 14532 27244
rect 14476 27134 14478 27186
rect 14530 27134 14532 27186
rect 14476 27122 14532 27134
rect 14700 27074 14756 28476
rect 14924 28532 14980 28542
rect 14924 28438 14980 28476
rect 15148 28418 15204 28430
rect 15148 28366 15150 28418
rect 15202 28366 15204 28418
rect 15148 27972 15204 28366
rect 15148 27906 15204 27916
rect 15372 28420 15428 28430
rect 14700 27022 14702 27074
rect 14754 27022 14756 27074
rect 14700 27010 14756 27022
rect 14812 27188 14868 27198
rect 14700 26516 14756 26526
rect 14812 26516 14868 27132
rect 15372 27074 15428 28364
rect 15596 28084 15652 29262
rect 15932 28868 15988 31836
rect 16044 31666 16100 31678
rect 16044 31614 16046 31666
rect 16098 31614 16100 31666
rect 16044 30996 16100 31614
rect 16156 31220 16212 31948
rect 16268 31220 16324 31230
rect 16212 31218 16324 31220
rect 16212 31166 16270 31218
rect 16322 31166 16324 31218
rect 16212 31164 16324 31166
rect 16156 31154 16212 31164
rect 16268 31154 16324 31164
rect 16044 30930 16100 30940
rect 16156 30994 16212 31006
rect 16156 30942 16158 30994
rect 16210 30942 16212 30994
rect 15708 28812 15988 28868
rect 16044 30548 16100 30558
rect 15708 28420 15764 28812
rect 15820 28644 15876 28654
rect 16044 28644 16100 30492
rect 16156 30212 16212 30942
rect 16268 30996 16324 31006
rect 16268 30770 16324 30940
rect 16268 30718 16270 30770
rect 16322 30718 16324 30770
rect 16268 30706 16324 30718
rect 16380 30548 16436 32844
rect 16492 32452 16548 32462
rect 16492 32358 16548 32396
rect 16604 32340 16660 32956
rect 16828 32564 16884 32574
rect 16828 32470 16884 32508
rect 16828 32340 16884 32350
rect 16604 32228 16660 32284
rect 16156 30146 16212 30156
rect 16268 30492 16436 30548
rect 16492 32172 16660 32228
rect 16716 32284 16828 32340
rect 16156 28644 16212 28654
rect 15820 28642 16212 28644
rect 15820 28590 15822 28642
rect 15874 28590 16158 28642
rect 16210 28590 16212 28642
rect 15820 28588 16212 28590
rect 15820 28578 15876 28588
rect 16156 28578 16212 28588
rect 16044 28420 16100 28430
rect 15708 28364 15988 28420
rect 15596 28018 15652 28028
rect 15484 27860 15540 27870
rect 15708 27860 15764 27870
rect 15484 27766 15540 27804
rect 15596 27858 15764 27860
rect 15596 27806 15710 27858
rect 15762 27806 15764 27858
rect 15596 27804 15764 27806
rect 15372 27022 15374 27074
rect 15426 27022 15428 27074
rect 15372 27010 15428 27022
rect 15148 26964 15204 27002
rect 15148 26898 15204 26908
rect 15260 26962 15316 26974
rect 15260 26910 15262 26962
rect 15314 26910 15316 26962
rect 15260 26908 15316 26910
rect 15596 26908 15652 27804
rect 15708 27794 15764 27804
rect 15820 27858 15876 27870
rect 15820 27806 15822 27858
rect 15874 27806 15876 27858
rect 15820 27636 15876 27806
rect 15820 27570 15876 27580
rect 15820 27300 15876 27310
rect 15932 27300 15988 28364
rect 15820 27298 15988 27300
rect 15820 27246 15822 27298
rect 15874 27246 15988 27298
rect 15820 27244 15988 27246
rect 15820 27234 15876 27244
rect 15708 27188 15764 27198
rect 15708 27076 15764 27132
rect 16044 27076 16100 28364
rect 16268 28196 16324 30492
rect 16492 30100 16548 32172
rect 16716 32004 16772 32284
rect 16828 32274 16884 32284
rect 16716 31938 16772 31948
rect 17052 32004 17108 32042
rect 17052 31938 17108 31948
rect 16604 31780 16660 31790
rect 17052 31780 17108 31790
rect 16604 31686 16660 31724
rect 16716 31778 17108 31780
rect 16716 31726 17054 31778
rect 17106 31726 17108 31778
rect 16716 31724 17108 31726
rect 16492 30034 16548 30044
rect 16716 29316 16772 31724
rect 17052 31714 17108 31724
rect 17052 31332 17108 31342
rect 17164 31332 17220 33068
rect 17108 31276 17220 31332
rect 17276 31332 17332 31342
rect 17052 31266 17108 31276
rect 16828 30996 16884 31006
rect 16828 30902 16884 30940
rect 17164 30884 17220 30894
rect 17276 30884 17332 31276
rect 17388 31106 17444 33516
rect 17500 33348 17556 33358
rect 17500 33254 17556 33292
rect 17612 32676 17668 33964
rect 17724 33908 17780 33918
rect 17780 33852 17892 33908
rect 17724 33842 17780 33852
rect 17388 31054 17390 31106
rect 17442 31054 17444 31106
rect 17388 31042 17444 31054
rect 17500 32620 17668 32676
rect 17276 30828 17444 30884
rect 17164 30322 17220 30828
rect 17164 30270 17166 30322
rect 17218 30270 17220 30322
rect 17164 30258 17220 30270
rect 15708 27074 16100 27076
rect 15708 27022 15710 27074
rect 15762 27022 16100 27074
rect 15708 27020 16100 27022
rect 16156 28140 16324 28196
rect 16380 29260 16772 29316
rect 17276 30100 17332 30110
rect 15708 27010 15764 27020
rect 14700 26514 14868 26516
rect 14700 26462 14702 26514
rect 14754 26462 14868 26514
rect 14700 26460 14868 26462
rect 15036 26852 15092 26862
rect 15260 26852 15652 26908
rect 15708 26852 15764 26862
rect 15036 26516 15092 26796
rect 15596 26740 15652 26750
rect 14700 26450 14756 26460
rect 15036 26422 15092 26460
rect 15260 26628 15316 26638
rect 14476 25844 14532 25854
rect 14476 25506 14532 25788
rect 14476 25454 14478 25506
rect 14530 25454 14532 25506
rect 14476 25442 14532 25454
rect 14700 25508 14756 25518
rect 14700 25394 14756 25452
rect 14700 25342 14702 25394
rect 14754 25342 14756 25394
rect 14700 25330 14756 25342
rect 15260 25282 15316 26572
rect 15372 26516 15428 26526
rect 15372 26402 15428 26460
rect 15596 26514 15652 26684
rect 15596 26462 15598 26514
rect 15650 26462 15652 26514
rect 15596 26450 15652 26462
rect 15708 26514 15764 26796
rect 15708 26462 15710 26514
rect 15762 26462 15764 26514
rect 15708 26450 15764 26462
rect 15820 26850 15876 26862
rect 15820 26798 15822 26850
rect 15874 26798 15876 26850
rect 15372 26350 15374 26402
rect 15426 26350 15428 26402
rect 15372 26338 15428 26350
rect 15708 26292 15764 26302
rect 15596 25506 15652 25518
rect 15596 25454 15598 25506
rect 15650 25454 15652 25506
rect 15596 25396 15652 25454
rect 15596 25330 15652 25340
rect 15260 25230 15262 25282
rect 15314 25230 15316 25282
rect 15260 25218 15316 25230
rect 14252 24770 14308 24780
rect 15708 24724 15764 26236
rect 15820 26290 15876 26798
rect 16156 26516 16212 28140
rect 16268 27634 16324 27646
rect 16268 27582 16270 27634
rect 16322 27582 16324 27634
rect 16268 27524 16324 27582
rect 16268 27458 16324 27468
rect 15820 26238 15822 26290
rect 15874 26238 15876 26290
rect 15820 25732 15876 26238
rect 15932 26460 16212 26516
rect 15932 25956 15988 26460
rect 16156 26404 16212 26460
rect 16156 26338 16212 26348
rect 16268 27300 16324 27310
rect 16044 26292 16100 26302
rect 16044 26198 16100 26236
rect 16268 25956 16324 27244
rect 16380 26852 16436 29260
rect 16716 28756 16772 28766
rect 16716 28532 16772 28700
rect 16716 28466 16772 28476
rect 16716 27972 16772 27982
rect 16772 27916 16884 27972
rect 16716 27878 16772 27916
rect 16604 27860 16660 27870
rect 16380 26786 16436 26796
rect 16492 27858 16660 27860
rect 16492 27806 16606 27858
rect 16658 27806 16660 27858
rect 16492 27804 16660 27806
rect 16492 26292 16548 27804
rect 16604 27794 16660 27804
rect 16716 27636 16772 27646
rect 16716 27542 16772 27580
rect 16828 27300 16884 27916
rect 17164 27300 17220 27310
rect 16828 27244 17164 27300
rect 17164 27186 17220 27244
rect 17164 27134 17166 27186
rect 17218 27134 17220 27186
rect 17164 27122 17220 27134
rect 16604 26852 16660 26862
rect 16604 26758 16660 26796
rect 16940 26852 16996 26862
rect 16492 26236 16772 26292
rect 15932 25890 15988 25900
rect 16156 25900 16324 25956
rect 16380 26180 16436 26190
rect 16156 25732 16212 25900
rect 15820 25666 15876 25676
rect 15932 25676 16212 25732
rect 16268 25732 16324 25742
rect 15932 24836 15988 25676
rect 16044 25508 16100 25518
rect 16044 25414 16100 25452
rect 16156 25396 16212 25406
rect 16044 24836 16100 24846
rect 15932 24834 16100 24836
rect 15932 24782 16046 24834
rect 16098 24782 16100 24834
rect 15932 24780 16100 24782
rect 15708 24668 15988 24724
rect 14028 23998 14030 24050
rect 14082 23998 14084 24050
rect 14028 23986 14084 23998
rect 14700 24276 14756 24286
rect 14700 23938 14756 24220
rect 15708 24164 15764 24174
rect 15148 24052 15204 24062
rect 15148 23958 15204 23996
rect 14700 23886 14702 23938
rect 14754 23886 14756 23938
rect 14700 23874 14756 23886
rect 15484 23940 15540 23950
rect 15148 23044 15204 23054
rect 15484 23044 15540 23884
rect 15708 23828 15764 24108
rect 15820 23828 15876 23838
rect 15708 23772 15820 23828
rect 15596 23380 15652 23390
rect 15708 23380 15764 23772
rect 15820 23762 15876 23772
rect 15596 23378 15764 23380
rect 15596 23326 15598 23378
rect 15650 23326 15764 23378
rect 15596 23324 15764 23326
rect 15932 23378 15988 24668
rect 15932 23326 15934 23378
rect 15986 23326 15988 23378
rect 15596 23314 15652 23324
rect 15820 23268 15876 23278
rect 15820 23174 15876 23212
rect 15148 23042 15540 23044
rect 15148 22990 15150 23042
rect 15202 22990 15540 23042
rect 15148 22988 15540 22990
rect 15148 22708 15204 22988
rect 15148 22642 15204 22652
rect 15596 22484 15652 22494
rect 15932 22484 15988 23326
rect 16044 22932 16100 24780
rect 16156 24050 16212 25340
rect 16268 25394 16324 25676
rect 16268 25342 16270 25394
rect 16322 25342 16324 25394
rect 16268 25330 16324 25342
rect 16380 24164 16436 26124
rect 16492 25620 16548 25630
rect 16716 25620 16772 26236
rect 16492 25618 16660 25620
rect 16492 25566 16494 25618
rect 16546 25566 16660 25618
rect 16492 25564 16660 25566
rect 16492 25554 16548 25564
rect 16492 24724 16548 24734
rect 16492 24630 16548 24668
rect 16380 24108 16548 24164
rect 16156 23998 16158 24050
rect 16210 23998 16212 24050
rect 16156 23986 16212 23998
rect 16380 23938 16436 23950
rect 16380 23886 16382 23938
rect 16434 23886 16436 23938
rect 16380 23492 16436 23886
rect 16156 23436 16436 23492
rect 16156 23378 16212 23436
rect 16156 23326 16158 23378
rect 16210 23326 16212 23378
rect 16156 23314 16212 23326
rect 16492 23380 16548 24108
rect 16604 23828 16660 25564
rect 16716 25554 16772 25564
rect 16828 26178 16884 26190
rect 16828 26126 16830 26178
rect 16882 26126 16884 26178
rect 16828 25508 16884 26126
rect 16940 26180 16996 26796
rect 16940 26114 16996 26124
rect 16716 24946 16772 24958
rect 16716 24894 16718 24946
rect 16770 24894 16772 24946
rect 16716 24724 16772 24894
rect 16716 24658 16772 24668
rect 16828 24612 16884 25452
rect 17276 24948 17332 30044
rect 17388 26908 17444 30828
rect 17500 30210 17556 32620
rect 17724 32564 17780 32574
rect 17724 32470 17780 32508
rect 17836 32340 17892 33852
rect 17948 33796 18004 34188
rect 18060 34178 18116 34188
rect 17948 33730 18004 33740
rect 18060 34020 18116 34030
rect 17948 33012 18004 33022
rect 17948 32564 18004 32956
rect 18060 32674 18116 33964
rect 18060 32622 18062 32674
rect 18114 32622 18116 32674
rect 18060 32610 18116 32622
rect 17948 32498 18004 32508
rect 18060 32452 18116 32462
rect 18060 32358 18116 32396
rect 17724 32284 17892 32340
rect 17612 31778 17668 31790
rect 17612 31726 17614 31778
rect 17666 31726 17668 31778
rect 17612 31332 17668 31726
rect 17724 31666 17780 32284
rect 18172 32116 18228 36092
rect 18284 34804 18340 36318
rect 18284 34738 18340 34748
rect 18396 36260 18452 36270
rect 18396 34356 18452 36204
rect 18508 35140 18564 36428
rect 18620 36260 18676 36270
rect 18620 35476 18676 36204
rect 18844 36036 18900 36876
rect 19292 36820 19348 44044
rect 19836 43932 20100 43942
rect 19892 43876 19940 43932
rect 19996 43876 20044 43932
rect 19836 43866 20100 43876
rect 19836 42364 20100 42374
rect 19892 42308 19940 42364
rect 19996 42308 20044 42364
rect 19836 42298 20100 42308
rect 20188 41972 20244 41982
rect 19964 41916 20188 41972
rect 19852 41858 19908 41870
rect 19852 41806 19854 41858
rect 19906 41806 19908 41858
rect 19516 41748 19572 41758
rect 19572 41692 19684 41748
rect 19516 41682 19572 41692
rect 19516 41188 19572 41198
rect 19516 40626 19572 41132
rect 19628 41186 19684 41692
rect 19852 41636 19908 41806
rect 19852 41570 19908 41580
rect 19628 41134 19630 41186
rect 19682 41134 19684 41186
rect 19628 41122 19684 41134
rect 19964 41186 20020 41916
rect 20188 41878 20244 41916
rect 19964 41134 19966 41186
rect 20018 41134 20020 41186
rect 19964 41122 20020 41134
rect 20188 41412 20244 41422
rect 19852 41076 19908 41086
rect 19852 40982 19908 41020
rect 19836 40796 20100 40806
rect 19892 40740 19940 40796
rect 19996 40740 20044 40796
rect 19836 40730 20100 40740
rect 19516 40574 19518 40626
rect 19570 40574 19572 40626
rect 19516 40562 19572 40574
rect 20188 40628 20244 41356
rect 20300 40964 20356 44716
rect 20412 42196 20468 47182
rect 20524 45444 20580 47404
rect 21308 46676 21364 56140
rect 21420 56130 21476 56140
rect 23324 56194 23380 56206
rect 23324 56142 23326 56194
rect 23378 56142 23380 56194
rect 23324 55636 23380 56142
rect 23548 56082 23604 56364
rect 25340 56364 25844 56420
rect 25340 56306 25396 56364
rect 25340 56254 25342 56306
rect 25394 56254 25396 56306
rect 25340 56242 25396 56254
rect 25564 56196 25620 56206
rect 23548 56030 23550 56082
rect 23602 56030 23604 56082
rect 23548 56018 23604 56030
rect 25452 56194 25620 56196
rect 25452 56142 25566 56194
rect 25618 56142 25620 56194
rect 25452 56140 25620 56142
rect 22988 55580 23380 55636
rect 21420 55300 21476 55310
rect 21420 55206 21476 55244
rect 22988 55298 23044 55580
rect 22988 55246 22990 55298
rect 23042 55246 23044 55298
rect 22988 55234 23044 55246
rect 23212 55412 23268 55422
rect 22876 55074 22932 55086
rect 22876 55022 22878 55074
rect 22930 55022 22932 55074
rect 22876 54516 22932 55022
rect 22764 54460 22876 54516
rect 21756 54402 21812 54414
rect 21756 54350 21758 54402
rect 21810 54350 21812 54402
rect 21756 53732 21812 54350
rect 21756 53666 21812 53676
rect 22428 53732 22484 53742
rect 22428 53638 22484 53676
rect 22652 53732 22708 53742
rect 22316 53620 22372 53630
rect 21980 53508 22036 53518
rect 21980 53414 22036 53452
rect 22316 52948 22372 53564
rect 22652 53508 22708 53676
rect 22652 53442 22708 53452
rect 22764 53060 22820 54460
rect 22876 54450 22932 54460
rect 22876 53844 22932 53854
rect 22876 53730 22932 53788
rect 22876 53678 22878 53730
rect 22930 53678 22932 53730
rect 22876 53666 22932 53678
rect 22764 52966 22820 53004
rect 22428 52948 22484 52958
rect 22316 52946 22484 52948
rect 22316 52894 22430 52946
rect 22482 52894 22484 52946
rect 22316 52892 22484 52894
rect 21756 52836 21812 52846
rect 21756 51490 21812 52780
rect 21756 51438 21758 51490
rect 21810 51438 21812 51490
rect 21756 51426 21812 51438
rect 22428 50820 22484 52892
rect 22988 52946 23044 52958
rect 22988 52894 22990 52946
rect 23042 52894 23044 52946
rect 22540 52836 22596 52846
rect 22540 52742 22596 52780
rect 21868 50596 21924 50606
rect 22092 50596 22148 50606
rect 21924 50594 22148 50596
rect 21924 50542 22094 50594
rect 22146 50542 22148 50594
rect 21924 50540 22148 50542
rect 21868 50502 21924 50540
rect 22092 50530 22148 50540
rect 22428 50482 22484 50764
rect 22988 50708 23044 52894
rect 22988 50642 23044 50652
rect 23100 52276 23156 52286
rect 22428 50430 22430 50482
rect 22482 50430 22484 50482
rect 22428 50418 22484 50430
rect 22204 49924 22260 49934
rect 21868 49028 21924 49038
rect 21868 48934 21924 48972
rect 22092 49026 22148 49038
rect 22092 48974 22094 49026
rect 22146 48974 22148 49026
rect 21868 48354 21924 48366
rect 21868 48302 21870 48354
rect 21922 48302 21924 48354
rect 21644 48244 21700 48254
rect 21644 47684 21700 48188
rect 21868 47908 21924 48302
rect 22092 48244 22148 48974
rect 22204 49026 22260 49868
rect 22652 49812 22708 49822
rect 23100 49812 23156 52220
rect 22652 49810 23156 49812
rect 22652 49758 22654 49810
rect 22706 49758 23102 49810
rect 23154 49758 23156 49810
rect 22652 49756 23156 49758
rect 22652 49746 22708 49756
rect 23100 49746 23156 49756
rect 23212 49588 23268 55356
rect 25340 55300 25396 55310
rect 25452 55300 25508 56140
rect 25564 56130 25620 56140
rect 25788 56082 25844 56364
rect 25788 56030 25790 56082
rect 25842 56030 25844 56082
rect 25788 56018 25844 56030
rect 27916 56306 27972 57148
rect 27916 56254 27918 56306
rect 27970 56254 27972 56306
rect 27916 56084 27972 56254
rect 29820 56420 29876 59200
rect 29820 56364 30324 56420
rect 29820 56306 29876 56364
rect 29820 56254 29822 56306
rect 29874 56254 29876 56306
rect 29820 56242 29876 56254
rect 27916 56018 27972 56028
rect 28364 56194 28420 56206
rect 28364 56142 28366 56194
rect 28418 56142 28420 56194
rect 28364 55468 28420 56142
rect 30044 56194 30100 56206
rect 30044 56142 30046 56194
rect 30098 56142 30100 56194
rect 28588 56084 28644 56094
rect 28588 55990 28644 56028
rect 30044 55468 30100 56142
rect 30268 56082 30324 56364
rect 31724 56308 31780 56318
rect 32060 56308 32116 59200
rect 34300 56308 34356 59200
rect 36540 56308 36596 59200
rect 38780 56642 38836 59200
rect 38780 56590 38782 56642
rect 38834 56590 38836 56642
rect 38780 56578 38836 56590
rect 39340 56642 39396 56654
rect 39340 56590 39342 56642
rect 39394 56590 39396 56642
rect 31724 56306 32340 56308
rect 31724 56254 31726 56306
rect 31778 56254 32340 56306
rect 31724 56252 32340 56254
rect 31724 56242 31780 56252
rect 32284 56194 32340 56252
rect 34300 56306 34580 56308
rect 34300 56254 34302 56306
rect 34354 56254 34580 56306
rect 34300 56252 34580 56254
rect 34300 56242 34356 56252
rect 32284 56142 32286 56194
rect 32338 56142 32340 56194
rect 32284 56130 32340 56142
rect 32620 56194 32676 56206
rect 32620 56142 32622 56194
rect 32674 56142 32676 56194
rect 30268 56030 30270 56082
rect 30322 56030 30324 56082
rect 30268 56018 30324 56030
rect 25340 55298 25508 55300
rect 25340 55246 25342 55298
rect 25394 55246 25508 55298
rect 25340 55244 25508 55246
rect 27692 55412 28420 55468
rect 29372 55412 30100 55468
rect 30492 55860 30548 55870
rect 27692 55298 27748 55412
rect 27692 55246 27694 55298
rect 27746 55246 27748 55298
rect 25340 55234 25396 55244
rect 27692 55234 27748 55246
rect 29260 55300 29316 55310
rect 29260 55206 29316 55244
rect 25228 55074 25284 55086
rect 25228 55022 25230 55074
rect 25282 55022 25284 55074
rect 23436 54516 23492 54526
rect 23436 53170 23492 54460
rect 23884 54402 23940 54414
rect 23884 54350 23886 54402
rect 23938 54350 23940 54402
rect 23660 53844 23716 53854
rect 23660 53750 23716 53788
rect 23772 53732 23828 53742
rect 23884 53732 23940 54350
rect 24892 54404 24948 54414
rect 23772 53730 24276 53732
rect 23772 53678 23774 53730
rect 23826 53678 24276 53730
rect 23772 53676 24276 53678
rect 23772 53666 23828 53676
rect 23436 53118 23438 53170
rect 23490 53118 23492 53170
rect 23436 53106 23492 53118
rect 23548 53506 23604 53518
rect 23548 53454 23550 53506
rect 23602 53454 23604 53506
rect 23548 52948 23604 53454
rect 23548 50484 23604 52892
rect 23996 53506 24052 53518
rect 23996 53454 23998 53506
rect 24050 53454 24052 53506
rect 23996 53060 24052 53454
rect 23884 51268 23940 51278
rect 23772 51266 23940 51268
rect 23772 51214 23886 51266
rect 23938 51214 23940 51266
rect 23772 51212 23940 51214
rect 23660 50708 23716 50718
rect 23660 50614 23716 50652
rect 23548 50418 23604 50428
rect 23772 50594 23828 51212
rect 23884 51202 23940 51212
rect 23772 50542 23774 50594
rect 23826 50542 23828 50594
rect 23772 49924 23828 50542
rect 23996 50482 24052 53004
rect 23996 50430 23998 50482
rect 24050 50430 24052 50482
rect 23996 50418 24052 50430
rect 24108 50596 24164 50606
rect 23772 49858 23828 49868
rect 22204 48974 22206 49026
rect 22258 48974 22260 49026
rect 22204 48962 22260 48974
rect 22988 49532 23268 49588
rect 24108 49698 24164 50540
rect 24220 50428 24276 53676
rect 24556 53730 24612 53742
rect 24556 53678 24558 53730
rect 24610 53678 24612 53730
rect 24556 53620 24612 53678
rect 24556 53554 24612 53564
rect 24892 53506 24948 54348
rect 25228 53844 25284 55022
rect 27580 55074 27636 55086
rect 27580 55022 27582 55074
rect 27634 55022 27636 55074
rect 25116 53788 25284 53844
rect 25340 54514 25396 54526
rect 25340 54462 25342 54514
rect 25394 54462 25396 54514
rect 24892 53454 24894 53506
rect 24946 53454 24948 53506
rect 24892 53442 24948 53454
rect 25004 53620 25060 53630
rect 25116 53620 25172 53788
rect 25004 53618 25172 53620
rect 25004 53566 25006 53618
rect 25058 53566 25172 53618
rect 25004 53564 25172 53566
rect 25228 53620 25284 53630
rect 25004 53508 25060 53564
rect 25228 53526 25284 53564
rect 24892 52612 24948 52622
rect 25004 52612 25060 53452
rect 24948 52556 25060 52612
rect 24892 52546 24948 52556
rect 25228 52164 25284 52174
rect 25228 52052 25284 52108
rect 25340 52052 25396 54462
rect 26012 54404 26068 54414
rect 26012 54310 26068 54348
rect 27580 54404 27636 55022
rect 29148 54740 29204 54750
rect 29148 54626 29204 54684
rect 29148 54574 29150 54626
rect 29202 54574 29204 54626
rect 28812 54516 28868 54526
rect 28812 54422 28868 54460
rect 26572 53844 26628 53854
rect 26348 53620 26404 53630
rect 26348 53526 26404 53564
rect 25676 53508 25732 53518
rect 25676 53414 25732 53452
rect 26236 53506 26292 53518
rect 26236 53454 26238 53506
rect 26290 53454 26292 53506
rect 25452 53060 25508 53070
rect 25452 52946 25508 53004
rect 25452 52894 25454 52946
rect 25506 52894 25508 52946
rect 25452 52882 25508 52894
rect 25900 52946 25956 52958
rect 25900 52894 25902 52946
rect 25954 52894 25956 52946
rect 25228 52050 25396 52052
rect 25228 51998 25230 52050
rect 25282 51998 25396 52050
rect 25228 51996 25396 51998
rect 25228 51986 25284 51996
rect 25340 51378 25396 51996
rect 25452 52500 25508 52510
rect 25452 52052 25508 52444
rect 25452 51986 25508 51996
rect 25340 51326 25342 51378
rect 25394 51326 25396 51378
rect 25340 51314 25396 51326
rect 25900 51268 25956 52894
rect 26124 52948 26180 52958
rect 26236 52948 26292 53454
rect 26460 53508 26516 53518
rect 26572 53508 26628 53788
rect 27580 53732 27636 54348
rect 28140 54402 28196 54414
rect 28140 54350 28142 54402
rect 28194 54350 28196 54402
rect 28140 53844 28196 54350
rect 29148 54292 29204 54574
rect 29148 53844 29204 54236
rect 29372 54180 29428 55412
rect 29932 55186 29988 55198
rect 29932 55134 29934 55186
rect 29986 55134 29988 55186
rect 29932 54738 29988 55134
rect 29932 54686 29934 54738
rect 29986 54686 29988 54738
rect 29932 54674 29988 54686
rect 29484 54626 29540 54638
rect 29484 54574 29486 54626
rect 29538 54574 29540 54626
rect 29484 54404 29540 54574
rect 29820 54514 29876 54526
rect 29820 54462 29822 54514
rect 29874 54462 29876 54514
rect 29820 54404 29876 54462
rect 30044 54516 30100 54526
rect 30044 54422 30100 54460
rect 29484 54348 29876 54404
rect 29372 54124 29764 54180
rect 29260 53844 29316 53854
rect 29148 53842 29316 53844
rect 29148 53790 29262 53842
rect 29314 53790 29316 53842
rect 29148 53788 29316 53790
rect 28140 53778 28196 53788
rect 29260 53778 29316 53788
rect 27580 53666 27636 53676
rect 26460 53506 26628 53508
rect 26460 53454 26462 53506
rect 26514 53454 26628 53506
rect 26460 53452 26628 53454
rect 26460 53442 26516 53452
rect 26180 52892 26292 52948
rect 26124 52854 26180 52892
rect 25900 51202 25956 51212
rect 26012 52834 26068 52846
rect 26012 52782 26014 52834
rect 26066 52782 26068 52834
rect 24444 50596 24500 50634
rect 24444 50530 24500 50540
rect 26012 50596 26068 52782
rect 26124 51268 26180 51278
rect 26124 51266 26516 51268
rect 26124 51214 26126 51266
rect 26178 51214 26516 51266
rect 26124 51212 26516 51214
rect 26124 51202 26180 51212
rect 26012 50530 26068 50540
rect 26236 50820 26292 50830
rect 26236 50594 26292 50764
rect 26460 50706 26516 51212
rect 26460 50654 26462 50706
rect 26514 50654 26516 50706
rect 26460 50642 26516 50654
rect 26236 50542 26238 50594
rect 26290 50542 26292 50594
rect 26236 50530 26292 50542
rect 24556 50484 24612 50494
rect 24780 50484 24836 50494
rect 24612 50482 24836 50484
rect 24612 50430 24782 50482
rect 24834 50430 24836 50482
rect 24612 50428 24836 50430
rect 26572 50428 26628 53452
rect 26684 53506 26740 53518
rect 26684 53454 26686 53506
rect 26738 53454 26740 53506
rect 26684 53060 26740 53454
rect 29260 53508 29316 53518
rect 29260 53170 29316 53452
rect 29260 53118 29262 53170
rect 29314 53118 29316 53170
rect 29260 53106 29316 53118
rect 26684 52966 26740 53004
rect 29708 53058 29764 54124
rect 29708 53006 29710 53058
rect 29762 53006 29764 53058
rect 29708 52994 29764 53006
rect 29820 53060 29876 54348
rect 30380 54290 30436 54302
rect 30380 54238 30382 54290
rect 30434 54238 30436 54290
rect 30380 53844 30436 54238
rect 30492 53956 30548 55804
rect 32060 55410 32116 55422
rect 32060 55358 32062 55410
rect 32114 55358 32116 55410
rect 31836 54628 31892 54638
rect 31892 54572 32004 54628
rect 31836 54534 31892 54572
rect 30604 54516 30660 54526
rect 30604 54514 31780 54516
rect 30604 54462 30606 54514
rect 30658 54462 31780 54514
rect 30604 54460 31780 54462
rect 30604 54450 30660 54460
rect 31724 54402 31780 54460
rect 31724 54350 31726 54402
rect 31778 54350 31780 54402
rect 31724 54338 31780 54350
rect 30492 53900 30660 53956
rect 30436 53788 30548 53844
rect 30380 53778 30436 53788
rect 30268 53508 30324 53518
rect 30044 53060 30100 53070
rect 29820 53004 30044 53060
rect 30044 52966 30100 53004
rect 30268 53058 30324 53452
rect 30268 53006 30270 53058
rect 30322 53006 30324 53058
rect 30268 52994 30324 53006
rect 27020 52946 27076 52958
rect 27020 52894 27022 52946
rect 27074 52894 27076 52946
rect 27020 52836 27076 52894
rect 30492 52946 30548 53788
rect 30492 52894 30494 52946
rect 30546 52894 30548 52946
rect 30492 52882 30548 52894
rect 27020 52770 27076 52780
rect 27468 52836 27524 52846
rect 27468 52742 27524 52780
rect 28476 52836 28532 52846
rect 27244 52276 27300 52286
rect 27244 52164 27300 52220
rect 27692 52164 27748 52174
rect 27244 52162 27748 52164
rect 27244 52110 27246 52162
rect 27298 52110 27694 52162
rect 27746 52110 27748 52162
rect 27244 52108 27748 52110
rect 27244 52098 27300 52108
rect 26796 52052 26852 52062
rect 26796 50820 26852 51996
rect 26684 50764 26796 50820
rect 26684 50594 26740 50764
rect 26796 50754 26852 50764
rect 26908 51380 26964 51390
rect 26684 50542 26686 50594
rect 26738 50542 26740 50594
rect 26684 50530 26740 50542
rect 26796 50596 26852 50606
rect 26796 50502 26852 50540
rect 24220 50372 24500 50428
rect 24556 50418 24612 50428
rect 24780 50418 24836 50428
rect 24108 49646 24110 49698
rect 24162 49646 24164 49698
rect 22540 48914 22596 48926
rect 22876 48916 22932 48926
rect 22540 48862 22542 48914
rect 22594 48862 22596 48914
rect 22428 48802 22484 48814
rect 22428 48750 22430 48802
rect 22482 48750 22484 48802
rect 22428 48356 22484 48750
rect 22428 48290 22484 48300
rect 22204 48244 22260 48254
rect 22092 48188 22204 48244
rect 22204 48178 22260 48188
rect 22428 48130 22484 48142
rect 22428 48078 22430 48130
rect 22482 48078 22484 48130
rect 22428 48020 22484 48078
rect 22428 47954 22484 47964
rect 21980 47908 22036 47918
rect 21868 47852 21980 47908
rect 21980 47842 22036 47852
rect 22540 47908 22596 48862
rect 22540 47684 22596 47852
rect 22764 48914 22932 48916
rect 22764 48862 22878 48914
rect 22930 48862 22932 48914
rect 22764 48860 22932 48862
rect 22764 48242 22820 48860
rect 22876 48850 22932 48860
rect 22988 48914 23044 49532
rect 22988 48862 22990 48914
rect 23042 48862 23044 48914
rect 22988 48850 23044 48862
rect 23212 48802 23268 48814
rect 23212 48750 23214 48802
rect 23266 48750 23268 48802
rect 22876 48692 22932 48702
rect 22876 48466 22932 48636
rect 22876 48414 22878 48466
rect 22930 48414 22932 48466
rect 22876 48402 22932 48414
rect 23212 48468 23268 48750
rect 23212 48402 23268 48412
rect 23884 48468 23940 48478
rect 23436 48354 23492 48366
rect 23436 48302 23438 48354
rect 23490 48302 23492 48354
rect 22764 48190 22766 48242
rect 22818 48190 22820 48242
rect 22764 47684 22820 48190
rect 22876 48244 22932 48254
rect 23100 48244 23156 48254
rect 23324 48244 23380 48254
rect 22932 48188 23044 48244
rect 22876 48178 22932 48188
rect 21644 47628 22260 47684
rect 21084 45780 21140 45790
rect 20636 45668 20692 45678
rect 20636 45666 20916 45668
rect 20636 45614 20638 45666
rect 20690 45614 20916 45666
rect 20636 45612 20916 45614
rect 20636 45602 20692 45612
rect 20524 45388 20692 45444
rect 20524 44882 20580 44894
rect 20524 44830 20526 44882
rect 20578 44830 20580 44882
rect 20524 44436 20580 44830
rect 20524 44370 20580 44380
rect 20636 43538 20692 45388
rect 20748 45332 20804 45342
rect 20748 45106 20804 45276
rect 20748 45054 20750 45106
rect 20802 45054 20804 45106
rect 20748 45042 20804 45054
rect 20860 44996 20916 45612
rect 20860 44930 20916 44940
rect 20972 44882 21028 44894
rect 20972 44830 20974 44882
rect 21026 44830 21028 44882
rect 20972 44548 21028 44830
rect 20972 44482 21028 44492
rect 20636 43486 20638 43538
rect 20690 43486 20692 43538
rect 20636 43474 20692 43486
rect 20748 44324 20804 44334
rect 21084 44324 21140 45724
rect 20748 42530 20804 44268
rect 20748 42478 20750 42530
rect 20802 42478 20804 42530
rect 20748 42420 20804 42478
rect 20748 42354 20804 42364
rect 20860 44268 21140 44324
rect 21196 45444 21252 45454
rect 20412 42140 20804 42196
rect 20412 41970 20468 41982
rect 20412 41918 20414 41970
rect 20466 41918 20468 41970
rect 20412 41076 20468 41918
rect 20636 41970 20692 41982
rect 20636 41918 20638 41970
rect 20690 41918 20692 41970
rect 20636 41636 20692 41918
rect 20636 41570 20692 41580
rect 20524 41076 20580 41086
rect 20412 41020 20524 41076
rect 20524 40982 20580 41020
rect 20300 40908 20468 40964
rect 20188 40562 20244 40572
rect 19516 39956 19572 39966
rect 19404 39396 19460 39406
rect 19404 39058 19460 39340
rect 19404 39006 19406 39058
rect 19458 39006 19460 39058
rect 19404 38994 19460 39006
rect 19516 39394 19572 39900
rect 20076 39844 20132 39854
rect 20076 39730 20132 39788
rect 20076 39678 20078 39730
rect 20130 39678 20132 39730
rect 20076 39666 20132 39678
rect 19516 39342 19518 39394
rect 19570 39342 19572 39394
rect 19516 38948 19572 39342
rect 20188 39396 20244 39406
rect 19836 39228 20100 39238
rect 19892 39172 19940 39228
rect 19996 39172 20044 39228
rect 19836 39162 20100 39172
rect 19516 38892 19684 38948
rect 19628 38276 19684 38892
rect 19740 38276 19796 38286
rect 19628 38220 19740 38276
rect 19628 38162 19684 38220
rect 19740 38210 19796 38220
rect 19628 38110 19630 38162
rect 19682 38110 19684 38162
rect 19628 38098 19684 38110
rect 19964 38052 20020 38062
rect 19964 37958 20020 37996
rect 19740 37940 19796 37950
rect 19740 37846 19796 37884
rect 19628 37828 19684 37838
rect 19404 37492 19460 37502
rect 19404 37398 19460 37436
rect 19068 36764 19348 36820
rect 19404 36932 19460 36942
rect 18956 36260 19012 36270
rect 18956 36166 19012 36204
rect 18844 35980 19012 36036
rect 18844 35812 18900 35822
rect 18620 35410 18676 35420
rect 18732 35698 18788 35710
rect 18732 35646 18734 35698
rect 18786 35646 18788 35698
rect 18508 35074 18564 35084
rect 18732 35026 18788 35646
rect 18844 35252 18900 35756
rect 18844 35186 18900 35196
rect 18732 34974 18734 35026
rect 18786 34974 18788 35026
rect 18732 34962 18788 34974
rect 18284 34300 18452 34356
rect 18508 34916 18564 34926
rect 18508 34354 18564 34860
rect 18844 34804 18900 34814
rect 18844 34710 18900 34748
rect 18956 34580 19012 35980
rect 19068 35922 19124 36764
rect 19180 36596 19236 36606
rect 19180 36372 19236 36540
rect 19292 36596 19348 36606
rect 19404 36596 19460 36876
rect 19292 36594 19460 36596
rect 19292 36542 19294 36594
rect 19346 36542 19460 36594
rect 19292 36540 19460 36542
rect 19292 36530 19348 36540
rect 19180 36316 19460 36372
rect 19068 35870 19070 35922
rect 19122 35870 19124 35922
rect 19068 35858 19124 35870
rect 19180 36148 19236 36158
rect 19180 35252 19236 36092
rect 19292 35812 19348 35822
rect 19292 35718 19348 35756
rect 19068 34692 19124 34702
rect 19068 34598 19124 34636
rect 18508 34302 18510 34354
rect 18562 34302 18564 34354
rect 18284 33460 18340 34300
rect 18508 34290 18564 34302
rect 18844 34524 19012 34580
rect 18396 34130 18452 34142
rect 18396 34078 18398 34130
rect 18450 34078 18452 34130
rect 18396 33908 18452 34078
rect 18396 33842 18452 33852
rect 18620 34130 18676 34142
rect 18620 34078 18622 34130
rect 18674 34078 18676 34130
rect 18284 33394 18340 33404
rect 18396 33346 18452 33358
rect 18396 33294 18398 33346
rect 18450 33294 18452 33346
rect 18284 33236 18340 33274
rect 18284 33170 18340 33180
rect 18284 33012 18340 33022
rect 18284 32228 18340 32956
rect 18396 32788 18452 33294
rect 18620 33124 18676 34078
rect 18844 33572 18900 34524
rect 19068 34132 19124 34142
rect 18956 33572 19012 33582
rect 18844 33570 19012 33572
rect 18844 33518 18958 33570
rect 19010 33518 19012 33570
rect 18844 33516 19012 33518
rect 18956 33506 19012 33516
rect 19068 33572 19124 34076
rect 19180 34020 19236 35196
rect 19404 35140 19460 36316
rect 19628 35924 19684 37772
rect 19836 37660 20100 37670
rect 19892 37604 19940 37660
rect 19996 37604 20044 37660
rect 19836 37594 20100 37604
rect 20076 37268 20132 37278
rect 20188 37268 20244 39340
rect 20300 38722 20356 38734
rect 20300 38670 20302 38722
rect 20354 38670 20356 38722
rect 20300 38500 20356 38670
rect 20412 38668 20468 40908
rect 20636 40962 20692 40974
rect 20636 40910 20638 40962
rect 20690 40910 20692 40962
rect 20636 40180 20692 40910
rect 20748 40964 20804 42140
rect 20860 41970 20916 44268
rect 21196 44100 21252 45388
rect 21308 44322 21364 46620
rect 21756 46564 21812 46574
rect 21812 46508 22036 46564
rect 21420 45892 21476 45902
rect 21644 45892 21700 45902
rect 21476 45890 21700 45892
rect 21476 45838 21646 45890
rect 21698 45838 21700 45890
rect 21476 45836 21700 45838
rect 21420 45826 21476 45836
rect 21644 45826 21700 45836
rect 21420 45666 21476 45678
rect 21420 45614 21422 45666
rect 21474 45614 21476 45666
rect 21420 45556 21476 45614
rect 21420 45490 21476 45500
rect 21532 45666 21588 45678
rect 21532 45614 21534 45666
rect 21586 45614 21588 45666
rect 21420 45332 21476 45342
rect 21532 45332 21588 45614
rect 21420 45330 21588 45332
rect 21420 45278 21422 45330
rect 21474 45278 21588 45330
rect 21420 45276 21588 45278
rect 21420 45266 21476 45276
rect 21644 45220 21700 45230
rect 21756 45220 21812 46508
rect 21980 45890 22036 46508
rect 22204 46002 22260 47628
rect 22204 45950 22206 46002
rect 22258 45950 22260 46002
rect 22204 45938 22260 45950
rect 22316 47628 22820 47684
rect 21980 45838 21982 45890
rect 22034 45838 22036 45890
rect 21980 45826 22036 45838
rect 21644 45218 21812 45220
rect 21644 45166 21646 45218
rect 21698 45166 21812 45218
rect 21644 45164 21812 45166
rect 21644 45154 21700 45164
rect 21308 44270 21310 44322
rect 21362 44270 21364 44322
rect 21308 44258 21364 44270
rect 21644 44660 21700 44670
rect 21644 44322 21700 44604
rect 21756 44548 21812 45164
rect 21756 44482 21812 44492
rect 21868 45106 21924 45118
rect 21868 45054 21870 45106
rect 21922 45054 21924 45106
rect 21644 44270 21646 44322
rect 21698 44270 21700 44322
rect 21644 44258 21700 44270
rect 21532 44210 21588 44222
rect 21532 44158 21534 44210
rect 21586 44158 21588 44210
rect 21532 44100 21588 44158
rect 21868 44212 21924 45054
rect 22316 45106 22372 47628
rect 22540 46900 22596 46910
rect 22316 45054 22318 45106
rect 22370 45054 22372 45106
rect 22316 45042 22372 45054
rect 22428 45666 22484 45678
rect 22428 45614 22430 45666
rect 22482 45614 22484 45666
rect 22092 44884 22148 44894
rect 21868 44146 21924 44156
rect 21980 44882 22148 44884
rect 21980 44830 22094 44882
rect 22146 44830 22148 44882
rect 21980 44828 22148 44830
rect 21196 44044 21588 44100
rect 21084 42868 21140 42878
rect 21532 42868 21588 44044
rect 21756 43650 21812 43662
rect 21756 43598 21758 43650
rect 21810 43598 21812 43650
rect 21756 43316 21812 43598
rect 21756 43250 21812 43260
rect 21756 42868 21812 42878
rect 21532 42866 21812 42868
rect 21532 42814 21758 42866
rect 21810 42814 21812 42866
rect 21532 42812 21812 42814
rect 20860 41918 20862 41970
rect 20914 41918 20916 41970
rect 20860 41636 20916 41918
rect 20972 41972 21028 41982
rect 20972 41878 21028 41916
rect 20860 41570 20916 41580
rect 20860 41412 20916 41422
rect 20860 41186 20916 41356
rect 20860 41134 20862 41186
rect 20914 41134 20916 41186
rect 20860 41122 20916 41134
rect 21084 41076 21140 42812
rect 21308 42532 21364 42542
rect 21308 42438 21364 42476
rect 21532 41860 21588 41870
rect 21532 41766 21588 41804
rect 21756 41636 21812 42812
rect 21980 41972 22036 44828
rect 22092 44818 22148 44828
rect 22092 44548 22148 44558
rect 22092 44454 22148 44492
rect 22316 43764 22372 43774
rect 22316 43670 22372 43708
rect 21980 41906 22036 41916
rect 22092 41970 22148 41982
rect 22092 41918 22094 41970
rect 22146 41918 22148 41970
rect 21868 41858 21924 41870
rect 21868 41806 21870 41858
rect 21922 41806 21924 41858
rect 21868 41748 21924 41806
rect 21980 41748 22036 41758
rect 21868 41692 21980 41748
rect 21980 41682 22036 41692
rect 21756 41580 21924 41636
rect 21756 41412 21812 41422
rect 21756 41318 21812 41356
rect 21420 41188 21476 41198
rect 21420 41094 21476 41132
rect 21532 41186 21588 41198
rect 21868 41188 21924 41580
rect 21532 41134 21534 41186
rect 21586 41134 21588 41186
rect 21084 41020 21364 41076
rect 20748 40908 21252 40964
rect 21084 40628 21140 40638
rect 21084 40534 21140 40572
rect 20636 39060 20692 40124
rect 21196 39396 21252 40908
rect 21308 39844 21364 41020
rect 21308 39618 21364 39788
rect 21532 39620 21588 41134
rect 21308 39566 21310 39618
rect 21362 39566 21364 39618
rect 21308 39554 21364 39566
rect 21420 39564 21588 39620
rect 21644 41132 21924 41188
rect 21980 41524 22036 41534
rect 21980 41186 22036 41468
rect 22092 41410 22148 41918
rect 22204 41970 22260 41982
rect 22204 41918 22206 41970
rect 22258 41918 22260 41970
rect 22204 41860 22260 41918
rect 22428 41970 22484 45614
rect 22540 45218 22596 46844
rect 22764 46562 22820 46574
rect 22764 46510 22766 46562
rect 22818 46510 22820 46562
rect 22652 46228 22708 46238
rect 22652 46002 22708 46172
rect 22652 45950 22654 46002
rect 22706 45950 22708 46002
rect 22652 45938 22708 45950
rect 22764 45556 22820 46510
rect 22764 45490 22820 45500
rect 22652 45332 22708 45342
rect 22652 45330 22932 45332
rect 22652 45278 22654 45330
rect 22706 45278 22932 45330
rect 22652 45276 22932 45278
rect 22652 45266 22708 45276
rect 22540 45166 22542 45218
rect 22594 45166 22596 45218
rect 22540 45154 22596 45166
rect 22876 45106 22932 45276
rect 22876 45054 22878 45106
rect 22930 45054 22932 45106
rect 22876 45042 22932 45054
rect 22988 45108 23044 48188
rect 23100 48242 23380 48244
rect 23100 48190 23102 48242
rect 23154 48190 23326 48242
rect 23378 48190 23380 48242
rect 23100 48188 23380 48190
rect 23100 48178 23156 48188
rect 23324 48178 23380 48188
rect 23436 48244 23492 48302
rect 23884 48354 23940 48412
rect 23884 48302 23886 48354
rect 23938 48302 23940 48354
rect 23884 48290 23940 48302
rect 23996 48354 24052 48366
rect 23996 48302 23998 48354
rect 24050 48302 24052 48354
rect 23436 48020 23492 48188
rect 23436 47954 23492 47964
rect 23660 48242 23716 48254
rect 23660 48190 23662 48242
rect 23714 48190 23716 48242
rect 23660 46116 23716 48190
rect 23996 48244 24052 48302
rect 23996 48178 24052 48188
rect 23996 48018 24052 48030
rect 23996 47966 23998 48018
rect 24050 47966 24052 48018
rect 23996 46900 24052 47966
rect 24108 47684 24164 49646
rect 24444 49140 24500 50372
rect 26460 50372 26628 50428
rect 25228 49924 25284 49934
rect 25228 49830 25284 49868
rect 25340 49586 25396 49598
rect 25340 49534 25342 49586
rect 25394 49534 25396 49586
rect 24556 49140 24612 49150
rect 24444 49138 24612 49140
rect 24444 49086 24558 49138
rect 24610 49086 24612 49138
rect 24444 49084 24612 49086
rect 24556 49074 24612 49084
rect 24668 49028 24724 49038
rect 24668 48934 24724 48972
rect 25340 48580 25396 49534
rect 25564 49028 25620 49038
rect 25564 48934 25620 48972
rect 26012 48914 26068 48926
rect 26012 48862 26014 48914
rect 26066 48862 26068 48914
rect 25340 48524 25956 48580
rect 25788 48356 25844 48366
rect 24556 48244 24612 48254
rect 24556 48150 24612 48188
rect 24108 47618 24164 47628
rect 24668 47236 24724 47246
rect 24668 47142 24724 47180
rect 25228 47236 25284 47246
rect 23996 46834 24052 46844
rect 24892 46900 24948 46910
rect 23660 46050 23716 46060
rect 24332 46562 24388 46574
rect 24780 46564 24836 46574
rect 24332 46510 24334 46562
rect 24386 46510 24388 46562
rect 23660 45778 23716 45790
rect 23660 45726 23662 45778
rect 23714 45726 23716 45778
rect 23100 45666 23156 45678
rect 23100 45614 23102 45666
rect 23154 45614 23156 45666
rect 23100 45444 23156 45614
rect 23100 45378 23156 45388
rect 23436 45332 23492 45342
rect 23436 45238 23492 45276
rect 23660 45220 23716 45726
rect 22988 45052 23380 45108
rect 23100 44882 23156 44894
rect 23100 44830 23102 44882
rect 23154 44830 23156 44882
rect 22988 44660 23044 44670
rect 22988 44322 23044 44604
rect 22988 44270 22990 44322
rect 23042 44270 23044 44322
rect 22988 44258 23044 44270
rect 22652 44212 22708 44222
rect 22652 44118 22708 44156
rect 23100 44100 23156 44830
rect 23100 44034 23156 44044
rect 23100 43428 23156 43438
rect 23100 43334 23156 43372
rect 22428 41918 22430 41970
rect 22482 41918 22484 41970
rect 22428 41906 22484 41918
rect 22652 42978 22708 42990
rect 22652 42926 22654 42978
rect 22706 42926 22708 42978
rect 22652 42530 22708 42926
rect 23212 42868 23268 42878
rect 22652 42478 22654 42530
rect 22706 42478 22708 42530
rect 22204 41794 22260 41804
rect 22092 41358 22094 41410
rect 22146 41358 22148 41410
rect 22092 41346 22148 41358
rect 21980 41134 21982 41186
rect 22034 41134 22036 41186
rect 21196 39340 21364 39396
rect 20636 39004 21028 39060
rect 20860 38836 20916 38846
rect 20636 38780 20860 38836
rect 20412 38612 20580 38668
rect 20300 38444 20468 38500
rect 20076 37266 20244 37268
rect 20076 37214 20078 37266
rect 20130 37214 20244 37266
rect 20076 37212 20244 37214
rect 20300 38050 20356 38062
rect 20300 37998 20302 38050
rect 20354 37998 20356 38050
rect 20076 37202 20132 37212
rect 19852 36596 19908 36606
rect 19852 36502 19908 36540
rect 20300 36484 20356 37998
rect 20412 36932 20468 38444
rect 20412 36866 20468 36876
rect 20412 36484 20468 36494
rect 20300 36482 20468 36484
rect 20300 36430 20414 36482
rect 20466 36430 20468 36482
rect 20300 36428 20468 36430
rect 20412 36418 20468 36428
rect 20300 36260 20356 36270
rect 20188 36204 20300 36260
rect 19836 36092 20100 36102
rect 19892 36036 19940 36092
rect 19996 36036 20044 36092
rect 19836 36026 20100 36036
rect 19740 35924 19796 35934
rect 19628 35922 19796 35924
rect 19628 35870 19742 35922
rect 19794 35870 19796 35922
rect 19628 35868 19796 35870
rect 19740 35858 19796 35868
rect 19852 35924 19908 35934
rect 19852 35308 19908 35868
rect 19404 35074 19460 35084
rect 19740 35252 19908 35308
rect 19964 35810 20020 35822
rect 19964 35758 19966 35810
rect 20018 35758 20020 35810
rect 19964 35364 20020 35758
rect 20076 35698 20132 35710
rect 20076 35646 20078 35698
rect 20130 35646 20132 35698
rect 20076 35588 20132 35646
rect 20076 35522 20132 35532
rect 19964 35298 20020 35308
rect 19404 34914 19460 34926
rect 19404 34862 19406 34914
rect 19458 34862 19460 34914
rect 19292 34690 19348 34702
rect 19292 34638 19294 34690
rect 19346 34638 19348 34690
rect 19292 34468 19348 34638
rect 19292 34402 19348 34412
rect 19180 33954 19236 33964
rect 19292 34132 19348 34142
rect 19068 33506 19124 33516
rect 19180 33460 19236 33470
rect 19068 33348 19124 33358
rect 18620 33058 18676 33068
rect 18844 33346 19124 33348
rect 18844 33294 19070 33346
rect 19122 33294 19124 33346
rect 18844 33292 19124 33294
rect 18396 32732 18564 32788
rect 18284 32172 18452 32228
rect 18172 32060 18340 32116
rect 17724 31614 17726 31666
rect 17778 31614 17780 31666
rect 17724 31444 17780 31614
rect 17724 31378 17780 31388
rect 17836 31668 17892 31678
rect 17612 31266 17668 31276
rect 17836 31218 17892 31612
rect 18060 31556 18116 31566
rect 17836 31166 17838 31218
rect 17890 31166 17892 31218
rect 17836 31154 17892 31166
rect 17948 31554 18116 31556
rect 17948 31502 18062 31554
rect 18114 31502 18116 31554
rect 17948 31500 18116 31502
rect 17612 31108 17668 31118
rect 17612 31014 17668 31052
rect 17836 30996 17892 31006
rect 17500 30158 17502 30210
rect 17554 30158 17556 30210
rect 17500 28756 17556 30158
rect 17724 30212 17780 30222
rect 17724 30118 17780 30156
rect 17500 28690 17556 28700
rect 17500 27860 17556 27870
rect 17500 27186 17556 27804
rect 17500 27134 17502 27186
rect 17554 27134 17556 27186
rect 17500 27122 17556 27134
rect 17724 27858 17780 27870
rect 17724 27806 17726 27858
rect 17778 27806 17780 27858
rect 17612 27076 17668 27086
rect 17388 26852 17556 26908
rect 17388 26290 17444 26302
rect 17388 26238 17390 26290
rect 17442 26238 17444 26290
rect 17388 26180 17444 26238
rect 17388 25506 17444 26124
rect 17388 25454 17390 25506
rect 17442 25454 17444 25506
rect 17388 25442 17444 25454
rect 17500 26068 17556 26852
rect 17612 26852 17668 27020
rect 17612 26786 17668 26796
rect 17724 26514 17780 27806
rect 17836 27860 17892 30940
rect 17948 30548 18004 31500
rect 18060 31490 18116 31500
rect 18172 31556 18228 31566
rect 18060 31220 18116 31258
rect 18060 31154 18116 31164
rect 18060 30996 18116 31006
rect 18172 30996 18228 31500
rect 18060 30994 18228 30996
rect 18060 30942 18062 30994
rect 18114 30942 18228 30994
rect 18060 30940 18228 30942
rect 18060 30930 18116 30940
rect 17948 30482 18004 30492
rect 18172 29876 18228 29886
rect 18172 28754 18228 29820
rect 18172 28702 18174 28754
rect 18226 28702 18228 28754
rect 18172 28420 18228 28702
rect 18284 28644 18340 32060
rect 18396 29876 18452 32172
rect 18508 31780 18564 32732
rect 18844 32562 18900 33292
rect 19068 33282 19124 33292
rect 18956 33124 19012 33134
rect 19180 33124 19236 33404
rect 18956 33030 19012 33068
rect 19068 33068 19236 33124
rect 19292 33348 19348 34076
rect 18844 32510 18846 32562
rect 18898 32510 18900 32562
rect 18844 32004 18900 32510
rect 18844 31938 18900 31948
rect 18508 31686 18564 31724
rect 18956 31554 19012 31566
rect 18956 31502 18958 31554
rect 19010 31502 19012 31554
rect 18508 31444 18564 31454
rect 18508 31106 18564 31388
rect 18956 31444 19012 31502
rect 18956 31378 19012 31388
rect 18732 31220 18788 31230
rect 18732 31126 18788 31164
rect 19068 31220 19124 33068
rect 19180 32788 19236 32798
rect 19292 32788 19348 33292
rect 19180 32786 19348 32788
rect 19180 32734 19182 32786
rect 19234 32734 19348 32786
rect 19180 32732 19348 32734
rect 19180 32722 19236 32732
rect 19068 31126 19124 31164
rect 19180 32116 19236 32126
rect 18508 31054 18510 31106
rect 18562 31054 18564 31106
rect 18508 31042 18564 31054
rect 18844 31108 18900 31118
rect 18844 31014 18900 31052
rect 18956 30996 19012 31006
rect 19180 30996 19236 32060
rect 18956 30902 19012 30940
rect 19068 30940 19236 30996
rect 19292 31444 19348 31454
rect 18956 29876 19012 29886
rect 18452 29820 18676 29876
rect 18396 29810 18452 29820
rect 18620 28980 18676 29820
rect 18956 29650 19012 29820
rect 18956 29598 18958 29650
rect 19010 29598 19012 29650
rect 18956 29586 19012 29598
rect 19068 29764 19124 30940
rect 19292 30884 19348 31388
rect 19292 30818 19348 30828
rect 19292 30660 19348 30670
rect 19068 29204 19124 29708
rect 19068 29138 19124 29148
rect 19180 30604 19292 30660
rect 19180 29986 19236 30604
rect 19292 30594 19348 30604
rect 19404 30100 19460 34862
rect 19740 34692 19796 35252
rect 20188 34916 20244 36204
rect 20300 36166 20356 36204
rect 20524 36036 20580 38612
rect 20636 38274 20692 38780
rect 20860 38770 20916 38780
rect 20636 38222 20638 38274
rect 20690 38222 20692 38274
rect 20636 38210 20692 38222
rect 20972 38722 21028 39004
rect 21308 38946 21364 39340
rect 21308 38894 21310 38946
rect 21362 38894 21364 38946
rect 21308 38882 21364 38894
rect 20972 38670 20974 38722
rect 21026 38670 21028 38722
rect 20748 36932 20804 36942
rect 20748 36482 20804 36876
rect 20748 36430 20750 36482
rect 20802 36430 20804 36482
rect 20748 36418 20804 36430
rect 20860 36484 20916 36494
rect 20412 35980 20580 36036
rect 20636 36258 20692 36270
rect 20636 36206 20638 36258
rect 20690 36206 20692 36258
rect 20300 35364 20356 35374
rect 20300 35026 20356 35308
rect 20300 34974 20302 35026
rect 20354 34974 20356 35026
rect 20300 34962 20356 34974
rect 20076 34860 20244 34916
rect 20412 34916 20468 35980
rect 20524 35810 20580 35822
rect 20524 35758 20526 35810
rect 20578 35758 20580 35810
rect 20524 35028 20580 35758
rect 20636 35700 20692 36206
rect 20860 35924 20916 36428
rect 20972 36036 21028 38670
rect 21196 38834 21252 38846
rect 21196 38782 21198 38834
rect 21250 38782 21252 38834
rect 21196 38668 21252 38782
rect 21196 38612 21364 38668
rect 21084 37604 21140 37614
rect 21084 37156 21140 37548
rect 21196 37378 21252 37390
rect 21196 37326 21198 37378
rect 21250 37326 21252 37378
rect 21196 37268 21252 37326
rect 21196 37202 21252 37212
rect 21084 37090 21140 37100
rect 20972 35970 21028 35980
rect 20860 35830 20916 35868
rect 20972 35700 21028 35710
rect 20636 35698 21028 35700
rect 20636 35646 20974 35698
rect 21026 35646 21028 35698
rect 20636 35644 21028 35646
rect 20860 35476 20916 35486
rect 20524 34972 20692 35028
rect 20412 34860 20580 34916
rect 20076 34692 20132 34860
rect 20188 34692 20244 34702
rect 20076 34690 20244 34692
rect 20076 34638 20190 34690
rect 20242 34638 20244 34690
rect 20076 34636 20244 34638
rect 19740 34626 19796 34636
rect 19836 34524 20100 34534
rect 19892 34468 19940 34524
rect 19996 34468 20044 34524
rect 19836 34458 20100 34468
rect 19964 34242 20020 34254
rect 19964 34190 19966 34242
rect 20018 34190 20020 34242
rect 19516 34132 19572 34142
rect 19516 34038 19572 34076
rect 19516 33124 19572 33134
rect 19516 33030 19572 33068
rect 19964 33124 20020 34190
rect 19964 33058 20020 33068
rect 19836 32956 20100 32966
rect 19892 32900 19940 32956
rect 19996 32900 20044 32956
rect 19836 32890 20100 32900
rect 20188 32900 20244 34636
rect 20412 34690 20468 34702
rect 20412 34638 20414 34690
rect 20466 34638 20468 34690
rect 20300 34130 20356 34142
rect 20300 34078 20302 34130
rect 20354 34078 20356 34130
rect 20300 34020 20356 34078
rect 20300 33458 20356 33964
rect 20300 33406 20302 33458
rect 20354 33406 20356 33458
rect 20300 33012 20356 33406
rect 20300 32946 20356 32956
rect 20188 32834 20244 32844
rect 19516 32676 19572 32686
rect 20412 32676 20468 34638
rect 19516 31778 19572 32620
rect 19852 32620 20468 32676
rect 19852 32450 19908 32620
rect 19852 32398 19854 32450
rect 19906 32398 19908 32450
rect 19852 32116 19908 32398
rect 19852 32050 19908 32060
rect 19964 32452 20020 32462
rect 19516 31726 19518 31778
rect 19570 31726 19572 31778
rect 19516 31668 19572 31726
rect 19516 31602 19572 31612
rect 19740 31556 19796 31566
rect 19964 31556 20020 32396
rect 20524 32004 20580 34860
rect 20412 31948 20580 32004
rect 20636 33236 20692 34972
rect 20860 34914 20916 35420
rect 20972 35364 21028 35644
rect 20972 35298 21028 35308
rect 20860 34862 20862 34914
rect 20914 34862 20916 34914
rect 20860 34850 20916 34862
rect 20972 34468 21028 34478
rect 20972 34132 21028 34412
rect 20972 34038 21028 34076
rect 21196 34130 21252 34142
rect 21196 34078 21198 34130
rect 21250 34078 21252 34130
rect 21196 33796 21252 34078
rect 21308 34132 21364 38612
rect 21420 37492 21476 39564
rect 21532 38836 21588 38846
rect 21532 38742 21588 38780
rect 21420 37426 21476 37436
rect 21532 37826 21588 37838
rect 21532 37774 21534 37826
rect 21586 37774 21588 37826
rect 21420 37156 21476 37166
rect 21420 37062 21476 37100
rect 21532 37044 21588 37774
rect 21532 36978 21588 36988
rect 21644 36596 21700 41132
rect 21980 40628 22036 41134
rect 22540 41076 22596 41086
rect 22540 40964 22596 41020
rect 21980 40562 22036 40572
rect 22428 40962 22596 40964
rect 22428 40910 22542 40962
rect 22594 40910 22596 40962
rect 22428 40908 22596 40910
rect 22316 40516 22372 40526
rect 22428 40516 22484 40908
rect 22540 40898 22596 40908
rect 22372 40460 22484 40516
rect 22316 40450 22372 40460
rect 22540 40404 22596 40414
rect 22540 40310 22596 40348
rect 22652 40180 22708 42478
rect 23100 42532 23156 42542
rect 22876 42196 22932 42206
rect 22876 41970 22932 42140
rect 22876 41918 22878 41970
rect 22930 41918 22932 41970
rect 22876 41906 22932 41918
rect 23100 41412 23156 42476
rect 23212 42532 23268 42812
rect 23324 42644 23380 45052
rect 23436 44434 23492 44446
rect 23436 44382 23438 44434
rect 23490 44382 23492 44434
rect 23436 44324 23492 44382
rect 23436 44258 23492 44268
rect 23660 44212 23716 45164
rect 24220 45780 24276 45790
rect 24332 45780 24388 46510
rect 24668 46562 24836 46564
rect 24668 46510 24782 46562
rect 24834 46510 24836 46562
rect 24668 46508 24836 46510
rect 24220 45778 24388 45780
rect 24220 45726 24222 45778
rect 24274 45726 24388 45778
rect 24220 45724 24388 45726
rect 24444 45890 24500 45902
rect 24444 45838 24446 45890
rect 24498 45838 24500 45890
rect 24220 44660 24276 45724
rect 24332 44996 24388 45006
rect 24332 44902 24388 44940
rect 24332 44660 24388 44670
rect 24220 44604 24332 44660
rect 23660 44146 23716 44156
rect 24220 44212 24276 44222
rect 24220 44118 24276 44156
rect 23772 43876 23828 43886
rect 23772 43762 23828 43820
rect 23772 43710 23774 43762
rect 23826 43710 23828 43762
rect 23772 43698 23828 43710
rect 23548 43652 23604 43662
rect 23436 43538 23492 43550
rect 23436 43486 23438 43538
rect 23490 43486 23492 43538
rect 23436 42978 23492 43486
rect 23436 42926 23438 42978
rect 23490 42926 23492 42978
rect 23436 42914 23492 42926
rect 23548 42868 23604 43596
rect 23996 43652 24052 43662
rect 23996 42978 24052 43596
rect 24220 43540 24276 43550
rect 24220 43316 24276 43484
rect 23996 42926 23998 42978
rect 24050 42926 24052 42978
rect 23996 42914 24052 42926
rect 24108 43092 24164 43102
rect 23660 42868 23716 42878
rect 23548 42866 23716 42868
rect 23548 42814 23662 42866
rect 23714 42814 23716 42866
rect 23548 42812 23716 42814
rect 23324 42588 23604 42644
rect 23212 42530 23380 42532
rect 23212 42478 23214 42530
rect 23266 42478 23380 42530
rect 23212 42476 23380 42478
rect 23212 42466 23268 42476
rect 22988 40964 23044 40974
rect 23100 40964 23156 41356
rect 22988 40962 23156 40964
rect 22988 40910 22990 40962
rect 23042 40910 23156 40962
rect 22988 40908 23156 40910
rect 23212 41858 23268 41870
rect 23212 41806 23214 41858
rect 23266 41806 23268 41858
rect 23212 41636 23268 41806
rect 22988 40898 23044 40908
rect 23212 40628 23268 41580
rect 23324 41860 23380 42476
rect 23324 41186 23380 41804
rect 23324 41134 23326 41186
rect 23378 41134 23380 41186
rect 23324 41076 23380 41134
rect 23324 41010 23380 41020
rect 23436 41748 23492 41758
rect 23212 40562 23268 40572
rect 23436 40404 23492 41692
rect 23436 40338 23492 40348
rect 22652 40114 22708 40124
rect 22204 39844 22260 39854
rect 22092 39730 22148 39742
rect 22092 39678 22094 39730
rect 22146 39678 22148 39730
rect 22092 38948 22148 39678
rect 22204 39058 22260 39788
rect 23324 39618 23380 39630
rect 23324 39566 23326 39618
rect 23378 39566 23380 39618
rect 22988 39396 23044 39406
rect 23324 39396 23380 39566
rect 22988 39394 23380 39396
rect 22988 39342 22990 39394
rect 23042 39342 23380 39394
rect 22988 39340 23380 39342
rect 22988 39330 23044 39340
rect 22204 39006 22206 39058
rect 22258 39006 22260 39058
rect 22204 38994 22260 39006
rect 21980 38836 22036 38846
rect 21980 38742 22036 38780
rect 21980 38276 22036 38286
rect 21980 37826 22036 38220
rect 21980 37774 21982 37826
rect 22034 37774 22036 37826
rect 21980 37604 22036 37774
rect 21980 37538 22036 37548
rect 21980 37380 22036 37390
rect 21868 36596 21924 36606
rect 21644 36540 21868 36596
rect 21532 36260 21588 36270
rect 21532 36258 21700 36260
rect 21532 36206 21534 36258
rect 21586 36206 21700 36258
rect 21532 36204 21700 36206
rect 21532 36194 21588 36204
rect 21420 35588 21476 35598
rect 21644 35588 21700 36204
rect 21476 35532 21588 35588
rect 21420 35522 21476 35532
rect 21532 34354 21588 35532
rect 21532 34302 21534 34354
rect 21586 34302 21588 34354
rect 21532 34290 21588 34302
rect 21644 34802 21700 35532
rect 21644 34750 21646 34802
rect 21698 34750 21700 34802
rect 21308 34066 21364 34076
rect 21196 33730 21252 33740
rect 20076 31892 20132 31902
rect 20076 31778 20132 31836
rect 20076 31726 20078 31778
rect 20130 31726 20132 31778
rect 20076 31714 20132 31726
rect 20188 31780 20244 31790
rect 20188 31686 20244 31724
rect 19180 29934 19182 29986
rect 19234 29934 19236 29986
rect 19180 28980 19236 29934
rect 18284 28588 18564 28644
rect 18396 28420 18452 28430
rect 18172 28354 18228 28364
rect 18284 28418 18452 28420
rect 18284 28366 18398 28418
rect 18450 28366 18452 28418
rect 18284 28364 18452 28366
rect 18172 28084 18228 28094
rect 18284 28084 18340 28364
rect 18396 28354 18452 28364
rect 18508 28196 18564 28588
rect 18620 28530 18676 28924
rect 19068 28924 19236 28980
rect 19292 30044 19460 30100
rect 19628 31554 20020 31556
rect 19628 31502 19742 31554
rect 19794 31502 20020 31554
rect 19628 31500 20020 31502
rect 20300 31556 20356 31566
rect 19628 30882 19684 31500
rect 19740 31490 19796 31500
rect 20300 31462 20356 31500
rect 19836 31388 20100 31398
rect 19892 31332 19940 31388
rect 19996 31332 20044 31388
rect 20412 31332 20468 31948
rect 19836 31322 20100 31332
rect 20188 31276 20468 31332
rect 20524 31780 20580 31790
rect 20636 31780 20692 33180
rect 20860 33684 20916 33694
rect 20748 33124 20804 33134
rect 20860 33124 20916 33628
rect 21644 33684 21700 34750
rect 21868 36258 21924 36540
rect 21868 36206 21870 36258
rect 21922 36206 21924 36258
rect 21868 34580 21924 36206
rect 21868 34514 21924 34524
rect 21980 34242 22036 37324
rect 22092 35700 22148 38892
rect 22652 38724 22708 38734
rect 22540 37826 22596 37838
rect 22540 37774 22542 37826
rect 22594 37774 22596 37826
rect 22540 37268 22596 37774
rect 22540 36482 22596 37212
rect 22652 37266 22708 38668
rect 22764 38722 22820 38734
rect 22764 38670 22766 38722
rect 22818 38670 22820 38722
rect 22764 37604 22820 38670
rect 22876 38388 22932 38398
rect 22876 38164 22932 38332
rect 22876 38070 22932 38108
rect 22764 37380 22820 37548
rect 22764 37314 22820 37324
rect 22652 37214 22654 37266
rect 22706 37214 22708 37266
rect 22652 37202 22708 37214
rect 22876 37266 22932 37278
rect 22876 37214 22878 37266
rect 22930 37214 22932 37266
rect 22540 36430 22542 36482
rect 22594 36430 22596 36482
rect 22540 36148 22596 36430
rect 22876 36148 22932 37214
rect 22988 37044 23044 37054
rect 22988 36370 23044 36988
rect 22988 36318 22990 36370
rect 23042 36318 23044 36370
rect 22988 36306 23044 36318
rect 22540 36082 22596 36092
rect 22764 36092 22932 36148
rect 22764 35700 22820 36092
rect 22876 35924 22932 35934
rect 22876 35810 22932 35868
rect 22876 35758 22878 35810
rect 22930 35758 22932 35810
rect 22876 35746 22932 35758
rect 22092 35644 22820 35700
rect 22988 35698 23044 35710
rect 22988 35646 22990 35698
rect 23042 35646 23044 35698
rect 22652 34916 22708 35644
rect 22988 35588 23044 35646
rect 21980 34190 21982 34242
rect 22034 34190 22036 34242
rect 21868 34132 21924 34142
rect 21868 33684 21924 34076
rect 21644 33618 21700 33628
rect 21756 33628 21924 33684
rect 20748 33122 20860 33124
rect 20748 33070 20750 33122
rect 20802 33070 20860 33122
rect 20748 33068 20860 33070
rect 20748 33058 20804 33068
rect 20860 33030 20916 33068
rect 21644 33122 21700 33134
rect 21644 33070 21646 33122
rect 21698 33070 21700 33122
rect 21644 32788 21700 33070
rect 21644 32722 21700 32732
rect 20860 32676 20916 32686
rect 20524 31778 20692 31780
rect 20524 31726 20526 31778
rect 20578 31726 20692 31778
rect 20524 31724 20692 31726
rect 20748 32620 20860 32676
rect 19740 31220 19796 31230
rect 19796 31164 20132 31220
rect 19740 31154 19796 31164
rect 20076 31106 20132 31164
rect 20076 31054 20078 31106
rect 20130 31054 20132 31106
rect 20076 31042 20132 31054
rect 19628 30830 19630 30882
rect 19682 30830 19684 30882
rect 18732 28868 18788 28878
rect 18732 28642 18788 28812
rect 18732 28590 18734 28642
rect 18786 28590 18788 28642
rect 18732 28578 18788 28590
rect 18844 28644 18900 28654
rect 18620 28478 18622 28530
rect 18674 28478 18676 28530
rect 18620 28466 18676 28478
rect 18172 28082 18340 28084
rect 18172 28030 18174 28082
rect 18226 28030 18340 28082
rect 18172 28028 18340 28030
rect 18396 28140 18564 28196
rect 18396 28082 18452 28140
rect 18396 28030 18398 28082
rect 18450 28030 18452 28082
rect 18172 28018 18228 28028
rect 18396 28018 18452 28030
rect 17836 27794 17892 27804
rect 17948 27860 18004 27870
rect 17948 27858 18228 27860
rect 17948 27806 17950 27858
rect 18002 27806 18228 27858
rect 17948 27804 18228 27806
rect 17948 27794 18004 27804
rect 18060 27412 18116 27422
rect 18172 27412 18228 27804
rect 18396 27858 18452 27870
rect 18396 27806 18398 27858
rect 18450 27806 18452 27858
rect 18396 27636 18452 27806
rect 18396 27570 18452 27580
rect 18508 27860 18564 27870
rect 18172 27356 18452 27412
rect 17948 27188 18004 27198
rect 17948 26628 18004 27132
rect 18060 27076 18116 27356
rect 18396 27186 18452 27356
rect 18396 27134 18398 27186
rect 18450 27134 18452 27186
rect 18396 27122 18452 27134
rect 18172 27076 18228 27086
rect 18060 27020 18172 27076
rect 17948 26562 18004 26572
rect 17724 26462 17726 26514
rect 17778 26462 17780 26514
rect 17724 26450 17780 26462
rect 17612 26404 17668 26414
rect 17612 26310 17668 26348
rect 17836 26290 17892 26302
rect 17836 26238 17838 26290
rect 17890 26238 17892 26290
rect 17836 26068 17892 26238
rect 17500 26012 17892 26068
rect 17948 26292 18004 26302
rect 17388 25172 17444 25182
rect 17500 25172 17556 26012
rect 17444 25116 17556 25172
rect 17612 25844 17668 25854
rect 17388 25106 17444 25116
rect 17276 24882 17332 24892
rect 17612 24946 17668 25788
rect 17724 25620 17780 25630
rect 17948 25620 18004 26236
rect 17724 25618 18004 25620
rect 17724 25566 17726 25618
rect 17778 25566 18004 25618
rect 17724 25564 18004 25566
rect 18060 25618 18116 25630
rect 18060 25566 18062 25618
rect 18114 25566 18116 25618
rect 17724 25284 17780 25564
rect 17724 25218 17780 25228
rect 17612 24894 17614 24946
rect 17666 24894 17668 24946
rect 17612 24882 17668 24894
rect 17836 24724 17892 24734
rect 17836 24630 17892 24668
rect 16828 24546 16884 24556
rect 18060 23938 18116 25566
rect 18172 25508 18228 27020
rect 18508 27074 18564 27804
rect 18732 27858 18788 27870
rect 18732 27806 18734 27858
rect 18786 27806 18788 27858
rect 18732 27188 18788 27806
rect 18732 27122 18788 27132
rect 18508 27022 18510 27074
rect 18562 27022 18564 27074
rect 18508 27010 18564 27022
rect 18844 27074 18900 28588
rect 19068 27636 19124 28924
rect 19180 28756 19236 28766
rect 19180 28662 19236 28700
rect 19068 27570 19124 27580
rect 19292 27972 19348 30044
rect 19628 29876 19684 30830
rect 20188 30884 20244 31276
rect 20524 31220 20580 31724
rect 20300 31164 20580 31220
rect 20636 31556 20692 31566
rect 20300 31106 20356 31164
rect 20300 31054 20302 31106
rect 20354 31054 20356 31106
rect 20300 31042 20356 31054
rect 20636 30994 20692 31500
rect 20636 30942 20638 30994
rect 20690 30942 20692 30994
rect 20636 30930 20692 30942
rect 20188 30828 20468 30884
rect 20076 30772 20132 30782
rect 19964 30436 20020 30446
rect 19964 30100 20020 30380
rect 19964 30006 20020 30044
rect 20076 30210 20132 30716
rect 20076 30158 20078 30210
rect 20130 30158 20132 30210
rect 20076 29988 20132 30158
rect 20076 29922 20132 29932
rect 19404 29820 19684 29876
rect 19836 29820 20100 29830
rect 19404 29428 19460 29820
rect 19892 29764 19940 29820
rect 19996 29764 20044 29820
rect 19836 29754 20100 29764
rect 19516 29652 19572 29662
rect 19740 29652 19796 29662
rect 19516 29650 19740 29652
rect 19516 29598 19518 29650
rect 19570 29598 19740 29650
rect 19516 29596 19740 29598
rect 19516 29586 19572 29596
rect 19404 29372 19572 29428
rect 19292 27634 19348 27916
rect 19292 27582 19294 27634
rect 19346 27582 19348 27634
rect 19292 27570 19348 27582
rect 19404 27860 19460 27870
rect 19292 27188 19348 27198
rect 19404 27188 19460 27804
rect 19292 27186 19460 27188
rect 19292 27134 19294 27186
rect 19346 27134 19460 27186
rect 19292 27132 19460 27134
rect 19292 27122 19348 27132
rect 19516 27076 19572 29372
rect 19740 29426 19796 29596
rect 20076 29652 20132 29662
rect 20076 29558 20132 29596
rect 20412 29540 20468 30828
rect 20748 30436 20804 32620
rect 20860 32610 20916 32620
rect 21644 32562 21700 32574
rect 21644 32510 21646 32562
rect 21698 32510 21700 32562
rect 21420 32452 21476 32462
rect 21644 32452 21700 32510
rect 21476 32396 21700 32452
rect 21420 32358 21476 32396
rect 21084 32340 21140 32350
rect 21140 32284 21252 32340
rect 21084 32274 21140 32284
rect 20860 31892 20916 31902
rect 20860 31798 20916 31836
rect 20972 31220 21028 31230
rect 20972 31218 21140 31220
rect 20972 31166 20974 31218
rect 21026 31166 21140 31218
rect 20972 31164 21140 31166
rect 20972 31154 21028 31164
rect 21084 31106 21140 31164
rect 21084 31054 21086 31106
rect 21138 31054 21140 31106
rect 21084 31042 21140 31054
rect 20860 30772 20916 30782
rect 21084 30772 21140 30782
rect 20860 30770 21140 30772
rect 20860 30718 20862 30770
rect 20914 30718 21086 30770
rect 21138 30718 21140 30770
rect 20860 30716 21140 30718
rect 20860 30706 20916 30716
rect 20748 30380 20916 30436
rect 20412 29446 20468 29484
rect 20748 30212 20804 30222
rect 19740 29374 19742 29426
rect 19794 29374 19796 29426
rect 19740 29362 19796 29374
rect 19964 29426 20020 29438
rect 19964 29374 19966 29426
rect 20018 29374 20020 29426
rect 19964 28980 20020 29374
rect 20188 29426 20244 29438
rect 20188 29374 20190 29426
rect 20242 29374 20244 29426
rect 19964 28914 20020 28924
rect 20076 29204 20132 29214
rect 20076 28756 20132 29148
rect 20188 29092 20244 29374
rect 20244 29036 20468 29092
rect 20188 29026 20244 29036
rect 20076 28754 20356 28756
rect 20076 28702 20078 28754
rect 20130 28702 20356 28754
rect 20076 28700 20356 28702
rect 20076 28690 20132 28700
rect 20188 28420 20244 28430
rect 20300 28420 20356 28700
rect 20412 28642 20468 29036
rect 20412 28590 20414 28642
rect 20466 28590 20468 28642
rect 20412 28578 20468 28590
rect 20748 28642 20804 30156
rect 20748 28590 20750 28642
rect 20802 28590 20804 28642
rect 20748 28578 20804 28590
rect 20524 28420 20580 28430
rect 20300 28418 20580 28420
rect 20300 28366 20526 28418
rect 20578 28366 20580 28418
rect 20300 28364 20580 28366
rect 19836 28252 20100 28262
rect 19892 28196 19940 28252
rect 19996 28196 20044 28252
rect 19836 28186 20100 28196
rect 19964 27860 20020 27870
rect 19964 27766 20020 27804
rect 20188 27860 20244 28364
rect 20524 28354 20580 28364
rect 20524 27972 20580 27982
rect 20524 27878 20580 27916
rect 20412 27860 20468 27870
rect 20188 27858 20468 27860
rect 20188 27806 20414 27858
rect 20466 27806 20468 27858
rect 20188 27804 20468 27806
rect 20188 27524 20244 27804
rect 20412 27794 20468 27804
rect 20860 27636 20916 30380
rect 20972 30324 21028 30716
rect 21084 30706 21140 30716
rect 20972 30258 21028 30268
rect 21196 29764 21252 32284
rect 21420 31668 21476 31678
rect 21420 31332 21476 31612
rect 21420 31266 21476 31276
rect 21308 31108 21364 31118
rect 21308 31106 21588 31108
rect 21308 31054 21310 31106
rect 21362 31054 21588 31106
rect 21308 31052 21588 31054
rect 21308 31042 21364 31052
rect 21420 30882 21476 30894
rect 21420 30830 21422 30882
rect 21474 30830 21476 30882
rect 21420 30772 21476 30830
rect 21420 30706 21476 30716
rect 21420 30436 21476 30446
rect 21420 30342 21476 30380
rect 21532 30210 21588 31052
rect 21756 30212 21812 33628
rect 21868 32674 21924 32686
rect 21868 32622 21870 32674
rect 21922 32622 21924 32674
rect 21868 31780 21924 32622
rect 21868 31714 21924 31724
rect 21868 31556 21924 31566
rect 21980 31556 22036 34190
rect 22540 34860 22708 34916
rect 22764 35532 23044 35588
rect 22204 34132 22260 34142
rect 22092 34130 22260 34132
rect 22092 34078 22206 34130
rect 22258 34078 22260 34130
rect 22092 34076 22260 34078
rect 22092 33460 22148 34076
rect 22204 34066 22260 34076
rect 22540 33908 22596 34860
rect 22764 34804 22820 35532
rect 22652 34692 22708 34702
rect 22652 34130 22708 34636
rect 22764 34690 22820 34748
rect 22764 34638 22766 34690
rect 22818 34638 22820 34690
rect 22764 34626 22820 34638
rect 22876 35364 22932 35374
rect 22876 34914 22932 35308
rect 22876 34862 22878 34914
rect 22930 34862 22932 34914
rect 22652 34078 22654 34130
rect 22706 34078 22708 34130
rect 22652 34066 22708 34078
rect 22092 33394 22148 33404
rect 22204 33852 22596 33908
rect 22652 33908 22708 33918
rect 22092 33236 22148 33246
rect 22092 33122 22148 33180
rect 22092 33070 22094 33122
rect 22146 33070 22148 33122
rect 22092 32228 22148 33070
rect 22092 32162 22148 32172
rect 21924 31500 22036 31556
rect 21868 31490 21924 31500
rect 21532 30158 21534 30210
rect 21586 30158 21588 30210
rect 21532 30146 21588 30158
rect 21644 30210 21812 30212
rect 21644 30158 21758 30210
rect 21810 30158 21812 30210
rect 21644 30156 21812 30158
rect 21196 29698 21252 29708
rect 21308 30098 21364 30110
rect 21308 30046 21310 30098
rect 21362 30046 21364 30098
rect 21308 29652 21364 30046
rect 21644 29988 21700 30156
rect 21756 30146 21812 30156
rect 21868 30882 21924 30894
rect 21868 30830 21870 30882
rect 21922 30830 21924 30882
rect 21868 30770 21924 30830
rect 21868 30718 21870 30770
rect 21922 30718 21924 30770
rect 21308 29586 21364 29596
rect 21420 29932 21700 29988
rect 21084 29540 21140 29550
rect 20972 29428 21028 29438
rect 20972 29334 21028 29372
rect 20188 27186 20244 27468
rect 20188 27134 20190 27186
rect 20242 27134 20244 27186
rect 20188 27122 20244 27134
rect 20524 27580 20916 27636
rect 20972 27970 21028 27982
rect 20972 27918 20974 27970
rect 21026 27918 21028 27970
rect 18844 27022 18846 27074
rect 18898 27022 18900 27074
rect 18844 27010 18900 27022
rect 19404 27020 19572 27076
rect 18284 26964 18340 27002
rect 19404 26908 19460 27020
rect 18284 26898 18340 26908
rect 19180 26852 19460 26908
rect 20300 26852 20356 26862
rect 18508 26404 18564 26414
rect 18508 26310 18564 26348
rect 19068 26178 19124 26190
rect 19068 26126 19070 26178
rect 19122 26126 19124 26178
rect 18396 25508 18452 25518
rect 18172 25506 18452 25508
rect 18172 25454 18398 25506
rect 18450 25454 18452 25506
rect 18172 25452 18452 25454
rect 18060 23886 18062 23938
rect 18114 23886 18116 23938
rect 18060 23874 18116 23886
rect 16940 23828 16996 23838
rect 16604 23826 16996 23828
rect 16604 23774 16942 23826
rect 16994 23774 16996 23826
rect 16604 23772 16996 23774
rect 16940 23762 16996 23772
rect 18172 23828 18228 23838
rect 18172 23734 18228 23772
rect 16716 23380 16772 23390
rect 16492 23378 16772 23380
rect 16492 23326 16718 23378
rect 16770 23326 16772 23378
rect 16492 23324 16772 23326
rect 18396 23380 18452 25452
rect 18844 25508 18900 25518
rect 18844 25414 18900 25452
rect 18620 25284 18676 25294
rect 18620 25060 18676 25228
rect 19068 25284 19124 26126
rect 19180 26180 19236 26852
rect 19836 26684 20100 26694
rect 19892 26628 19940 26684
rect 19996 26628 20044 26684
rect 19836 26618 20100 26628
rect 19180 26114 19236 26124
rect 19852 26180 19908 26190
rect 19740 25620 19796 25630
rect 19740 25506 19796 25564
rect 19740 25454 19742 25506
rect 19794 25454 19796 25506
rect 19740 25442 19796 25454
rect 19852 25508 19908 26124
rect 20300 26178 20356 26796
rect 20300 26126 20302 26178
rect 20354 26126 20356 26178
rect 19964 25844 20020 25854
rect 19964 25618 20020 25788
rect 19964 25566 19966 25618
rect 20018 25566 20020 25618
rect 19964 25554 20020 25566
rect 20300 25620 20356 26126
rect 20300 25554 20356 25564
rect 19852 25442 19908 25452
rect 20076 25506 20132 25518
rect 20076 25454 20078 25506
rect 20130 25454 20132 25506
rect 19068 25218 19124 25228
rect 20076 25284 20132 25454
rect 20076 25218 20132 25228
rect 20412 25394 20468 25406
rect 20412 25342 20414 25394
rect 20466 25342 20468 25394
rect 19836 25116 20100 25126
rect 19892 25060 19940 25116
rect 19996 25060 20044 25116
rect 18620 25004 19236 25060
rect 19836 25050 20100 25060
rect 18508 24612 18564 24622
rect 18508 24518 18564 24556
rect 19068 24612 19124 24622
rect 18620 23380 18676 23390
rect 18396 23378 18676 23380
rect 18396 23326 18622 23378
rect 18674 23326 18676 23378
rect 18396 23324 18676 23326
rect 16716 23314 16772 23324
rect 18620 23314 18676 23324
rect 19068 23378 19124 24556
rect 19068 23326 19070 23378
rect 19122 23326 19124 23378
rect 19068 23314 19124 23326
rect 19180 23266 19236 25004
rect 19180 23214 19182 23266
rect 19234 23214 19236 23266
rect 19180 23202 19236 23214
rect 19292 24834 19348 24846
rect 20412 24836 20468 25342
rect 19292 24782 19294 24834
rect 19346 24782 19348 24834
rect 17612 23042 17668 23054
rect 17612 22990 17614 23042
rect 17666 22990 17668 23042
rect 16156 22932 16212 22942
rect 16044 22876 16156 22932
rect 16156 22866 16212 22876
rect 17612 22932 17668 22990
rect 17612 22866 17668 22876
rect 19068 22932 19124 22942
rect 19292 22932 19348 24782
rect 20300 24834 20468 24836
rect 20300 24782 20414 24834
rect 20466 24782 20468 24834
rect 20300 24780 20468 24782
rect 19964 24724 20020 24734
rect 19740 24052 19796 24062
rect 19740 23958 19796 23996
rect 19964 23938 20020 24668
rect 19964 23886 19966 23938
rect 20018 23886 20020 23938
rect 19964 23874 20020 23886
rect 20188 23940 20244 23950
rect 20188 23846 20244 23884
rect 20300 23938 20356 24780
rect 20412 24770 20468 24780
rect 20524 24052 20580 27580
rect 20972 26908 21028 27918
rect 20860 26852 21028 26908
rect 20748 26180 20804 26190
rect 20748 26086 20804 26124
rect 20748 24164 20804 24174
rect 20860 24164 20916 26852
rect 21084 26516 21140 29484
rect 21420 28866 21476 29932
rect 21532 29428 21588 29438
rect 21532 29334 21588 29372
rect 21420 28814 21422 28866
rect 21474 28814 21476 28866
rect 21420 28802 21476 28814
rect 21868 28868 21924 30718
rect 21980 30098 22036 30110
rect 21980 30046 21982 30098
rect 22034 30046 22036 30098
rect 21980 29652 22036 30046
rect 21980 29586 22036 29596
rect 21980 29428 22036 29438
rect 22036 29372 22148 29428
rect 21980 29334 22036 29372
rect 21868 28812 22036 28868
rect 21868 28642 21924 28654
rect 21868 28590 21870 28642
rect 21922 28590 21924 28642
rect 21532 28532 21588 28542
rect 21868 28532 21924 28590
rect 21588 28476 21924 28532
rect 21532 28438 21588 28476
rect 21084 26290 21140 26460
rect 21084 26238 21086 26290
rect 21138 26238 21140 26290
rect 21084 26226 21140 26238
rect 21420 28418 21476 28430
rect 21420 28366 21422 28418
rect 21474 28366 21476 28418
rect 21420 26964 21476 28366
rect 21644 27972 21700 27982
rect 21644 27878 21700 27916
rect 20748 24162 20916 24164
rect 20748 24110 20750 24162
rect 20802 24110 20916 24162
rect 20748 24108 20916 24110
rect 21084 24722 21140 24734
rect 21084 24670 21086 24722
rect 21138 24670 21140 24722
rect 20748 24098 20804 24108
rect 20524 23986 20580 23996
rect 20300 23886 20302 23938
rect 20354 23886 20356 23938
rect 20300 23874 20356 23886
rect 21084 23940 21140 24670
rect 21084 23828 21140 23884
rect 21308 23828 21364 23838
rect 21084 23826 21364 23828
rect 21084 23774 21310 23826
rect 21362 23774 21364 23826
rect 21084 23772 21364 23774
rect 21308 23762 21364 23772
rect 21084 23604 21140 23614
rect 19836 23548 20100 23558
rect 19892 23492 19940 23548
rect 19996 23492 20044 23548
rect 19836 23482 20100 23492
rect 21084 23378 21140 23548
rect 21084 23326 21086 23378
rect 21138 23326 21140 23378
rect 21084 23314 21140 23326
rect 21308 23268 21364 23278
rect 21420 23268 21476 26908
rect 21868 26850 21924 26862
rect 21868 26798 21870 26850
rect 21922 26798 21924 26850
rect 21644 26292 21700 26302
rect 21868 26292 21924 26798
rect 21700 26236 21924 26292
rect 21644 26198 21700 26236
rect 21980 26180 22036 28812
rect 22092 26292 22148 29372
rect 22092 26198 22148 26236
rect 21868 26124 22036 26180
rect 21756 25506 21812 25518
rect 21756 25454 21758 25506
rect 21810 25454 21812 25506
rect 21532 25284 21588 25294
rect 21756 25284 21812 25454
rect 21588 25228 21812 25284
rect 21532 25190 21588 25228
rect 21868 24050 21924 26124
rect 22092 24836 22148 24846
rect 22092 24742 22148 24780
rect 21868 23998 21870 24050
rect 21922 23998 21924 24050
rect 21868 23604 21924 23998
rect 22204 24724 22260 33852
rect 22316 33348 22372 33358
rect 22316 32674 22372 33292
rect 22316 32622 22318 32674
rect 22370 32622 22372 32674
rect 22316 32610 22372 32622
rect 22540 33122 22596 33134
rect 22540 33070 22542 33122
rect 22594 33070 22596 33122
rect 22540 32564 22596 33070
rect 22540 32498 22596 32508
rect 22316 31780 22372 31790
rect 22316 31686 22372 31724
rect 22540 31780 22596 31790
rect 22540 31220 22596 31724
rect 22652 31556 22708 33852
rect 22764 33012 22820 33022
rect 22764 32674 22820 32956
rect 22764 32622 22766 32674
rect 22818 32622 22820 32674
rect 22764 32610 22820 32622
rect 22764 31780 22820 31790
rect 22764 31686 22820 31724
rect 22876 31668 22932 34862
rect 22988 33460 23044 33470
rect 22988 33122 23044 33404
rect 22988 33070 22990 33122
rect 23042 33070 23044 33122
rect 22988 32564 23044 33070
rect 23100 32676 23156 39340
rect 23212 38724 23268 38734
rect 23212 38630 23268 38668
rect 23324 38612 23380 38622
rect 23324 38052 23380 38556
rect 23548 38052 23604 42588
rect 23660 42532 23716 42812
rect 23660 42466 23716 42476
rect 23884 42642 23940 42654
rect 23884 42590 23886 42642
rect 23938 42590 23940 42642
rect 23884 42420 23940 42590
rect 23996 42532 24052 42542
rect 23996 42438 24052 42476
rect 23884 42354 23940 42364
rect 23660 42308 23716 42318
rect 23660 42194 23716 42252
rect 23660 42142 23662 42194
rect 23714 42142 23716 42194
rect 23660 42130 23716 42142
rect 23884 41074 23940 41086
rect 23884 41022 23886 41074
rect 23938 41022 23940 41074
rect 23884 40516 23940 41022
rect 24108 40628 24164 43036
rect 23884 40450 23940 40460
rect 23996 40626 24164 40628
rect 23996 40574 24110 40626
rect 24162 40574 24164 40626
rect 23996 40572 24164 40574
rect 23884 39508 23940 39518
rect 23884 39414 23940 39452
rect 23772 38834 23828 38846
rect 23772 38782 23774 38834
rect 23826 38782 23828 38834
rect 23772 38668 23828 38782
rect 23996 38668 24052 40572
rect 24108 40562 24164 40572
rect 24220 42308 24276 43260
rect 24220 40068 24276 42252
rect 24332 41076 24388 44604
rect 24444 44324 24500 45838
rect 24556 45780 24612 45790
rect 24556 45686 24612 45724
rect 24668 45220 24724 46508
rect 24780 46498 24836 46508
rect 24668 45154 24724 45164
rect 24780 45890 24836 45902
rect 24780 45838 24782 45890
rect 24834 45838 24836 45890
rect 24668 44994 24724 45006
rect 24668 44942 24670 44994
rect 24722 44942 24724 44994
rect 24668 44660 24724 44942
rect 24668 44594 24724 44604
rect 24668 44436 24724 44446
rect 24668 44342 24724 44380
rect 24556 44324 24612 44334
rect 24444 44322 24556 44324
rect 24444 44270 24446 44322
rect 24498 44270 24556 44322
rect 24444 44268 24556 44270
rect 24444 44258 24500 44268
rect 24556 43876 24612 44268
rect 24556 43650 24612 43820
rect 24556 43598 24558 43650
rect 24610 43598 24612 43650
rect 24556 43586 24612 43598
rect 24668 43316 24724 43326
rect 24668 43222 24724 43260
rect 24780 43092 24836 45838
rect 24892 45778 24948 46844
rect 25228 46674 25284 47180
rect 25228 46622 25230 46674
rect 25282 46622 25284 46674
rect 25228 46610 25284 46622
rect 24892 45726 24894 45778
rect 24946 45726 24948 45778
rect 24892 45714 24948 45726
rect 25676 45332 25732 45342
rect 25452 45330 25732 45332
rect 25452 45278 25678 45330
rect 25730 45278 25732 45330
rect 25452 45276 25732 45278
rect 25004 44100 25060 44110
rect 24556 43036 24836 43092
rect 24892 44044 25004 44100
rect 24444 42756 24500 42766
rect 24444 42662 24500 42700
rect 24556 41298 24612 43036
rect 24668 42754 24724 42766
rect 24668 42702 24670 42754
rect 24722 42702 24724 42754
rect 24668 42420 24724 42702
rect 24668 42354 24724 42364
rect 24668 41860 24724 41870
rect 24892 41860 24948 44044
rect 25004 44006 25060 44044
rect 25340 43650 25396 43662
rect 25340 43598 25342 43650
rect 25394 43598 25396 43650
rect 25228 43428 25284 43438
rect 25004 43426 25284 43428
rect 25004 43374 25230 43426
rect 25282 43374 25284 43426
rect 25004 43372 25284 43374
rect 25004 42978 25060 43372
rect 25228 43362 25284 43372
rect 25004 42926 25006 42978
rect 25058 42926 25060 42978
rect 25004 42914 25060 42926
rect 25004 42756 25060 42766
rect 25060 42700 25172 42756
rect 25004 42690 25060 42700
rect 24668 41858 24948 41860
rect 24668 41806 24670 41858
rect 24722 41806 24948 41858
rect 24668 41804 24948 41806
rect 24668 41524 24724 41804
rect 24668 41458 24724 41468
rect 24556 41246 24558 41298
rect 24610 41246 24612 41298
rect 24556 41234 24612 41246
rect 24892 41412 24948 41422
rect 24892 41186 24948 41356
rect 24892 41134 24894 41186
rect 24946 41134 24948 41186
rect 24892 41122 24948 41134
rect 24332 41020 24836 41076
rect 23772 38612 24052 38668
rect 23996 38610 24052 38612
rect 23996 38558 23998 38610
rect 24050 38558 24052 38610
rect 23996 38546 24052 38558
rect 24108 40012 24276 40068
rect 24108 38276 24164 40012
rect 24668 39396 24724 39406
rect 24220 38948 24276 38958
rect 24220 38854 24276 38892
rect 24668 38834 24724 39340
rect 24668 38782 24670 38834
rect 24722 38782 24724 38834
rect 24556 38722 24612 38734
rect 24556 38670 24558 38722
rect 24610 38670 24612 38722
rect 24556 38668 24612 38670
rect 24108 38210 24164 38220
rect 24444 38612 24612 38668
rect 23548 37996 24052 38052
rect 23324 37986 23380 37996
rect 23436 37826 23492 37838
rect 23436 37774 23438 37826
rect 23490 37774 23492 37826
rect 23212 37266 23268 37278
rect 23212 37214 23214 37266
rect 23266 37214 23268 37266
rect 23212 36932 23268 37214
rect 23436 37268 23492 37774
rect 23772 37826 23828 37838
rect 23772 37774 23774 37826
rect 23826 37774 23828 37826
rect 23548 37268 23604 37278
rect 23436 37266 23604 37268
rect 23436 37214 23550 37266
rect 23602 37214 23604 37266
rect 23436 37212 23604 37214
rect 23212 36866 23268 36876
rect 23436 36932 23492 36942
rect 23436 35586 23492 36876
rect 23548 35924 23604 37212
rect 23548 35858 23604 35868
rect 23548 35700 23604 35710
rect 23548 35698 23716 35700
rect 23548 35646 23550 35698
rect 23602 35646 23716 35698
rect 23548 35644 23716 35646
rect 23548 35634 23604 35644
rect 23436 35534 23438 35586
rect 23490 35534 23492 35586
rect 23436 35522 23492 35534
rect 23548 34130 23604 34142
rect 23548 34078 23550 34130
rect 23602 34078 23604 34130
rect 23548 33572 23604 34078
rect 23436 33516 23604 33572
rect 23324 33460 23380 33470
rect 23324 33366 23380 33404
rect 23436 33348 23492 33516
rect 23660 33460 23716 35644
rect 23772 35252 23828 37774
rect 23884 36258 23940 36270
rect 23884 36206 23886 36258
rect 23938 36206 23940 36258
rect 23884 35810 23940 36206
rect 23884 35758 23886 35810
rect 23938 35758 23940 35810
rect 23884 35746 23940 35758
rect 23772 35186 23828 35196
rect 23884 35364 23940 35374
rect 23772 34916 23828 34926
rect 23884 34916 23940 35308
rect 23772 34914 23940 34916
rect 23772 34862 23774 34914
rect 23826 34862 23940 34914
rect 23772 34860 23940 34862
rect 23772 34580 23828 34860
rect 23772 33908 23828 34524
rect 23996 34354 24052 37996
rect 24108 38050 24164 38062
rect 24108 37998 24110 38050
rect 24162 37998 24164 38050
rect 24108 37828 24164 37998
rect 24220 37940 24276 37950
rect 24332 37940 24388 37950
rect 24220 37938 24332 37940
rect 24220 37886 24222 37938
rect 24274 37886 24332 37938
rect 24220 37884 24332 37886
rect 24220 37874 24276 37884
rect 24108 37762 24164 37772
rect 24220 36482 24276 36494
rect 24220 36430 24222 36482
rect 24274 36430 24276 36482
rect 24220 36372 24276 36430
rect 23996 34302 23998 34354
rect 24050 34302 24052 34354
rect 23996 34290 24052 34302
rect 24108 35028 24164 35038
rect 23772 33842 23828 33852
rect 23884 34242 23940 34254
rect 23884 34190 23886 34242
rect 23938 34190 23940 34242
rect 23436 33282 23492 33292
rect 23548 33404 23716 33460
rect 23212 33124 23268 33134
rect 23212 33030 23268 33068
rect 23436 33122 23492 33134
rect 23436 33070 23438 33122
rect 23490 33070 23492 33122
rect 23436 32788 23492 33070
rect 23436 32722 23492 32732
rect 23100 32610 23156 32620
rect 22988 31892 23044 32508
rect 22988 31826 23044 31836
rect 23436 32228 23492 32238
rect 23436 31890 23492 32172
rect 23436 31838 23438 31890
rect 23490 31838 23492 31890
rect 23436 31826 23492 31838
rect 23100 31668 23156 31678
rect 22876 31612 23044 31668
rect 22652 31500 22932 31556
rect 22316 31164 22596 31220
rect 22652 31332 22708 31342
rect 22316 28642 22372 31164
rect 22540 30210 22596 30222
rect 22540 30158 22542 30210
rect 22594 30158 22596 30210
rect 22540 30100 22596 30158
rect 22540 30034 22596 30044
rect 22652 30098 22708 31276
rect 22652 30046 22654 30098
rect 22706 30046 22708 30098
rect 22652 29876 22708 30046
rect 22652 29810 22708 29820
rect 22428 29540 22484 29550
rect 22428 29446 22484 29484
rect 22316 28590 22318 28642
rect 22370 28590 22372 28642
rect 22316 28578 22372 28590
rect 22876 28642 22932 31500
rect 22876 28590 22878 28642
rect 22930 28590 22932 28642
rect 22876 28532 22932 28590
rect 22876 28466 22932 28476
rect 22652 27748 22708 27758
rect 22652 26908 22708 27692
rect 22988 26908 23044 31612
rect 23100 29428 23156 31612
rect 23212 31332 23268 31342
rect 23548 31332 23604 33404
rect 23772 33348 23828 33358
rect 23884 33348 23940 34190
rect 23996 34132 24052 34142
rect 23996 34038 24052 34076
rect 23772 33346 23940 33348
rect 23772 33294 23774 33346
rect 23826 33294 23940 33346
rect 23772 33292 23940 33294
rect 23660 32562 23716 32574
rect 23660 32510 23662 32562
rect 23714 32510 23716 32562
rect 23660 31780 23716 32510
rect 23660 31714 23716 31724
rect 23212 30884 23268 31276
rect 23212 30818 23268 30828
rect 23324 31276 23604 31332
rect 23212 30100 23268 30110
rect 23212 30006 23268 30044
rect 23100 29362 23156 29372
rect 22540 26852 22708 26908
rect 22764 26852 23044 26908
rect 23324 26908 23380 31276
rect 23772 30996 23828 33292
rect 24108 31444 24164 34972
rect 24220 34802 24276 36316
rect 24332 35812 24388 37884
rect 24332 35746 24388 35756
rect 24220 34750 24222 34802
rect 24274 34750 24276 34802
rect 24220 33012 24276 34750
rect 24220 32946 24276 32956
rect 24444 33012 24500 38612
rect 24444 32946 24500 32956
rect 24556 37604 24612 37614
rect 24332 32004 24388 32014
rect 23884 31388 24164 31444
rect 24220 31666 24276 31678
rect 24220 31614 24222 31666
rect 24274 31614 24276 31666
rect 23884 31220 23940 31388
rect 24220 31332 24276 31614
rect 23884 31126 23940 31164
rect 24108 31276 24276 31332
rect 24108 30996 24164 31276
rect 23660 30940 24164 30996
rect 24220 30996 24276 31006
rect 23548 30212 23604 30222
rect 23548 29988 23604 30156
rect 23548 29922 23604 29932
rect 23436 29876 23492 29886
rect 23436 29652 23492 29820
rect 23548 29652 23604 29662
rect 23436 29650 23604 29652
rect 23436 29598 23550 29650
rect 23602 29598 23604 29650
rect 23436 29596 23604 29598
rect 23548 29586 23604 29596
rect 23436 28644 23492 28654
rect 23436 28530 23492 28588
rect 23436 28478 23438 28530
rect 23490 28478 23492 28530
rect 23436 28466 23492 28478
rect 23548 28642 23604 28654
rect 23548 28590 23550 28642
rect 23602 28590 23604 28642
rect 23548 27748 23604 28590
rect 23548 27682 23604 27692
rect 23660 26908 23716 30940
rect 24220 30902 24276 30940
rect 24332 30772 24388 31948
rect 24444 31780 24500 31790
rect 24444 31556 24500 31724
rect 24444 31490 24500 31500
rect 24444 31108 24500 31118
rect 24444 31014 24500 31052
rect 24556 30882 24612 37548
rect 24668 37380 24724 38782
rect 24668 37314 24724 37324
rect 24668 35028 24724 35038
rect 24668 34354 24724 34972
rect 24668 34302 24670 34354
rect 24722 34302 24724 34354
rect 24668 34290 24724 34302
rect 24668 32452 24724 32462
rect 24668 32358 24724 32396
rect 24556 30830 24558 30882
rect 24610 30830 24612 30882
rect 24556 30818 24612 30830
rect 24668 31106 24724 31118
rect 24668 31054 24670 31106
rect 24722 31054 24724 31106
rect 24220 30716 24388 30772
rect 24108 30100 24164 30110
rect 24108 30006 24164 30044
rect 23996 29986 24052 29998
rect 23996 29934 23998 29986
rect 24050 29934 24052 29986
rect 23884 29764 23940 29774
rect 23884 29650 23940 29708
rect 23884 29598 23886 29650
rect 23938 29598 23940 29650
rect 23884 29586 23940 29598
rect 23772 27188 23828 27198
rect 23772 27094 23828 27132
rect 23324 26852 23492 26908
rect 22428 25394 22484 25406
rect 22428 25342 22430 25394
rect 22482 25342 22484 25394
rect 21868 23538 21924 23548
rect 21980 23940 22036 23950
rect 22204 23940 22260 24668
rect 21980 23938 22260 23940
rect 21980 23886 21982 23938
rect 22034 23886 22260 23938
rect 21980 23884 22260 23886
rect 21644 23380 21700 23390
rect 21980 23380 22036 23884
rect 21644 23378 22036 23380
rect 21644 23326 21646 23378
rect 21698 23326 22036 23378
rect 21644 23324 22036 23326
rect 22204 23380 22260 23884
rect 22316 24724 22372 24734
rect 22428 24724 22484 25342
rect 22540 25284 22596 26852
rect 22652 26180 22708 26190
rect 22764 26180 22820 26852
rect 22652 26178 22820 26180
rect 22652 26126 22654 26178
rect 22706 26126 22820 26178
rect 22652 26124 22820 26126
rect 23100 26292 23156 26302
rect 23100 26178 23156 26236
rect 23100 26126 23102 26178
rect 23154 26126 23156 26178
rect 22652 25396 22708 26124
rect 22652 25330 22708 25340
rect 22764 25732 22820 25742
rect 22540 25218 22596 25228
rect 22764 24946 22820 25676
rect 23100 25172 23156 26126
rect 23100 25106 23156 25116
rect 23324 25844 23380 25854
rect 22764 24894 22766 24946
rect 22818 24894 22820 24946
rect 22764 24882 22820 24894
rect 22316 24722 22484 24724
rect 22316 24670 22318 24722
rect 22370 24670 22484 24722
rect 22316 24668 22484 24670
rect 22316 24164 22372 24668
rect 22316 23938 22372 24108
rect 23324 24050 23380 25788
rect 23436 25618 23492 26852
rect 23548 26852 23716 26908
rect 23548 25732 23604 26852
rect 23548 25666 23604 25676
rect 23436 25566 23438 25618
rect 23490 25566 23492 25618
rect 23436 25554 23492 25566
rect 23660 25508 23716 25518
rect 23660 25414 23716 25452
rect 23548 25396 23604 25406
rect 23548 25302 23604 25340
rect 23324 23998 23326 24050
rect 23378 23998 23380 24050
rect 23324 23986 23380 23998
rect 23772 24276 23828 24286
rect 22316 23886 22318 23938
rect 22370 23886 22372 23938
rect 22316 23874 22372 23886
rect 23772 23938 23828 24220
rect 23772 23886 23774 23938
rect 23826 23886 23828 23938
rect 23772 23874 23828 23886
rect 23996 23492 24052 29934
rect 24108 29652 24164 29662
rect 24108 29558 24164 29596
rect 24220 29428 24276 30716
rect 24556 30212 24612 30222
rect 24556 30098 24612 30156
rect 24556 30046 24558 30098
rect 24610 30046 24612 30098
rect 24556 30034 24612 30046
rect 24332 29764 24388 29774
rect 24332 29650 24388 29708
rect 24332 29598 24334 29650
rect 24386 29598 24388 29650
rect 24332 29586 24388 29598
rect 24108 29372 24276 29428
rect 24444 29426 24500 29438
rect 24444 29374 24446 29426
rect 24498 29374 24500 29426
rect 24108 28642 24164 29372
rect 24444 29316 24500 29374
rect 24444 29250 24500 29260
rect 24108 28590 24110 28642
rect 24162 28590 24164 28642
rect 24108 24612 24164 28590
rect 24220 28532 24276 28542
rect 24220 28438 24276 28476
rect 24332 28420 24388 28430
rect 24332 28326 24388 28364
rect 24668 28084 24724 31054
rect 24668 28018 24724 28028
rect 24668 27746 24724 27758
rect 24668 27694 24670 27746
rect 24722 27694 24724 27746
rect 24668 27636 24724 27694
rect 24668 27570 24724 27580
rect 24780 27298 24836 41020
rect 25116 41074 25172 42700
rect 25340 42084 25396 43598
rect 25452 43204 25508 45276
rect 25676 45266 25732 45276
rect 25564 45106 25620 45118
rect 25564 45054 25566 45106
rect 25618 45054 25620 45106
rect 25564 44996 25620 45054
rect 25564 43708 25620 44940
rect 25788 44884 25844 48300
rect 25900 47458 25956 48524
rect 25900 47406 25902 47458
rect 25954 47406 25956 47458
rect 25900 47394 25956 47406
rect 26012 48356 26068 48862
rect 26012 47346 26068 48300
rect 26460 48354 26516 50372
rect 26908 48804 26964 51324
rect 27580 51268 27636 51278
rect 27356 50708 27412 50718
rect 27356 50614 27412 50652
rect 27580 49922 27636 51212
rect 27692 50428 27748 52108
rect 28476 52052 28532 52780
rect 30156 52834 30212 52846
rect 30156 52782 30158 52834
rect 30210 52782 30212 52834
rect 29596 52722 29652 52734
rect 29596 52670 29598 52722
rect 29650 52670 29652 52722
rect 29372 52164 29428 52174
rect 29372 52070 29428 52108
rect 29596 52052 29652 52670
rect 30156 52274 30212 52782
rect 30156 52222 30158 52274
rect 30210 52222 30212 52274
rect 30156 52210 30212 52222
rect 28476 51996 28644 52052
rect 28252 51268 28308 51278
rect 28252 51174 28308 51212
rect 27692 50372 27972 50428
rect 27580 49870 27582 49922
rect 27634 49870 27636 49922
rect 27580 49858 27636 49870
rect 27692 49586 27748 49598
rect 27692 49534 27694 49586
rect 27746 49534 27748 49586
rect 27244 49026 27300 49038
rect 27244 48974 27246 49026
rect 27298 48974 27300 49026
rect 27132 48916 27188 48926
rect 26908 48748 27076 48804
rect 26460 48302 26462 48354
rect 26514 48302 26516 48354
rect 26460 48290 26516 48302
rect 26572 48244 26628 48254
rect 26572 48150 26628 48188
rect 26012 47294 26014 47346
rect 26066 47294 26068 47346
rect 25900 45220 25956 45230
rect 25900 45126 25956 45164
rect 25676 44828 25844 44884
rect 25676 44324 25732 44828
rect 25788 44548 25844 44558
rect 26012 44548 26068 47294
rect 26908 47236 26964 47246
rect 27020 47236 27076 48748
rect 27132 48802 27188 48860
rect 27132 48750 27134 48802
rect 27186 48750 27188 48802
rect 27132 48738 27188 48750
rect 26908 47234 27076 47236
rect 26908 47182 26910 47234
rect 26962 47182 27076 47234
rect 26908 47180 27076 47182
rect 27132 48242 27188 48254
rect 27132 48190 27134 48242
rect 27186 48190 27188 48242
rect 26908 47170 26964 47180
rect 27132 47068 27188 48190
rect 27020 47012 27188 47068
rect 26796 45892 26852 45902
rect 26796 45798 26852 45836
rect 26236 45218 26292 45230
rect 26236 45166 26238 45218
rect 26290 45166 26292 45218
rect 26124 45108 26180 45118
rect 26124 45014 26180 45052
rect 25788 44546 26068 44548
rect 25788 44494 25790 44546
rect 25842 44494 26068 44546
rect 25788 44492 26068 44494
rect 25788 44482 25844 44492
rect 26124 44436 26180 44446
rect 26124 44342 26180 44380
rect 25676 44268 25844 44324
rect 25564 43652 25732 43708
rect 25564 43538 25620 43550
rect 25564 43486 25566 43538
rect 25618 43486 25620 43538
rect 25564 43428 25620 43486
rect 25564 43362 25620 43372
rect 25452 43148 25620 43204
rect 25564 42756 25620 43148
rect 25564 42662 25620 42700
rect 25452 42644 25508 42654
rect 25452 42550 25508 42588
rect 25116 41022 25118 41074
rect 25170 41022 25172 41074
rect 25116 41010 25172 41022
rect 25228 42028 25396 42084
rect 25452 42420 25508 42430
rect 25676 42420 25732 43652
rect 25788 43538 25844 44268
rect 26236 44212 26292 45166
rect 26348 44660 26404 44670
rect 26348 44322 26404 44604
rect 27020 44436 27076 47012
rect 27132 45556 27188 45566
rect 27132 44546 27188 45500
rect 27132 44494 27134 44546
rect 27186 44494 27188 44546
rect 27132 44482 27188 44494
rect 27020 44370 27076 44380
rect 26348 44270 26350 44322
rect 26402 44270 26404 44322
rect 26348 44258 26404 44270
rect 26684 44324 26740 44334
rect 26684 44230 26740 44268
rect 25788 43486 25790 43538
rect 25842 43486 25844 43538
rect 25788 43474 25844 43486
rect 25900 44156 26292 44212
rect 26460 44212 26516 44222
rect 25508 42364 25732 42420
rect 25116 40628 25172 40638
rect 25116 40292 25172 40572
rect 25228 40514 25284 42028
rect 25340 41860 25396 41870
rect 25452 41860 25508 42364
rect 25340 41858 25508 41860
rect 25340 41806 25342 41858
rect 25394 41806 25508 41858
rect 25340 41804 25508 41806
rect 25340 41748 25396 41804
rect 25340 41682 25396 41692
rect 25228 40462 25230 40514
rect 25282 40462 25284 40514
rect 25228 40450 25284 40462
rect 25116 40236 25284 40292
rect 25004 39284 25060 39294
rect 25004 38668 25060 39228
rect 25116 39060 25172 39070
rect 25116 38966 25172 39004
rect 25228 38836 25284 40236
rect 25340 40178 25396 40190
rect 25340 40126 25342 40178
rect 25394 40126 25396 40178
rect 25340 39284 25396 40126
rect 25340 39218 25396 39228
rect 25564 40178 25620 40190
rect 25564 40126 25566 40178
rect 25618 40126 25620 40178
rect 25564 39284 25620 40126
rect 25564 39218 25620 39228
rect 25676 40180 25732 40190
rect 25228 38780 25396 38836
rect 24892 38612 25060 38668
rect 24892 37940 24948 38612
rect 24892 37874 24948 37884
rect 25004 38500 25060 38510
rect 25004 32002 25060 38444
rect 25228 37492 25284 37502
rect 25228 37398 25284 37436
rect 25228 37156 25284 37166
rect 25228 35698 25284 37100
rect 25340 36708 25396 38780
rect 25564 38724 25620 38762
rect 25564 38658 25620 38668
rect 25564 38164 25620 38174
rect 25452 37378 25508 37390
rect 25452 37326 25454 37378
rect 25506 37326 25508 37378
rect 25452 37268 25508 37326
rect 25452 37202 25508 37212
rect 25564 37378 25620 38108
rect 25676 37604 25732 40124
rect 25788 39396 25844 39406
rect 25788 38834 25844 39340
rect 25900 39060 25956 44156
rect 26348 43988 26404 43998
rect 26236 43932 26348 43988
rect 26236 43650 26292 43932
rect 26348 43922 26404 43932
rect 26236 43598 26238 43650
rect 26290 43598 26292 43650
rect 26236 43586 26292 43598
rect 26460 43540 26516 44156
rect 26572 43652 26628 43662
rect 26572 43558 26628 43596
rect 26348 43484 26516 43540
rect 26348 40516 26404 43484
rect 26796 42532 26852 42542
rect 26572 41860 26628 41870
rect 26572 41766 26628 41804
rect 26348 40450 26404 40460
rect 26460 41076 26516 41086
rect 26124 40290 26180 40302
rect 26124 40238 26126 40290
rect 26178 40238 26180 40290
rect 26124 40068 26180 40238
rect 26348 40180 26404 40190
rect 26348 40086 26404 40124
rect 25900 38994 25956 39004
rect 26012 40012 26124 40068
rect 25788 38782 25790 38834
rect 25842 38782 25844 38834
rect 25788 38724 25844 38782
rect 26012 38834 26068 40012
rect 26124 40002 26180 40012
rect 26460 39730 26516 41020
rect 26684 40628 26740 40638
rect 26796 40628 26852 42476
rect 27244 42196 27300 48974
rect 27356 48356 27412 48366
rect 27356 48354 27636 48356
rect 27356 48302 27358 48354
rect 27410 48302 27636 48354
rect 27356 48300 27636 48302
rect 27356 48290 27412 48300
rect 27356 47460 27412 47470
rect 27356 47366 27412 47404
rect 27356 45780 27412 45790
rect 27356 45686 27412 45724
rect 27580 45330 27636 48300
rect 27692 47460 27748 49534
rect 27692 47394 27748 47404
rect 27804 48914 27860 48926
rect 27804 48862 27806 48914
rect 27858 48862 27860 48914
rect 27804 46002 27860 48862
rect 27916 47012 27972 50372
rect 28588 48132 28644 51996
rect 29596 51986 29652 51996
rect 30492 51380 30548 51390
rect 30604 51380 30660 53900
rect 31948 53172 32004 54572
rect 32060 54290 32116 55358
rect 32620 55298 32676 56142
rect 34524 56194 34580 56252
rect 36540 56306 36820 56308
rect 36540 56254 36542 56306
rect 36594 56254 36820 56306
rect 36540 56252 36820 56254
rect 36540 56242 36596 56252
rect 34524 56142 34526 56194
rect 34578 56142 34580 56194
rect 34524 56130 34580 56142
rect 34860 56194 34916 56206
rect 34860 56142 34862 56194
rect 34914 56142 34916 56194
rect 32620 55246 32622 55298
rect 32674 55246 32676 55298
rect 32620 55234 32676 55246
rect 33180 55300 33236 55310
rect 33628 55300 33684 55310
rect 33180 55206 33236 55244
rect 33516 55244 33628 55300
rect 32620 55074 32676 55086
rect 32620 55022 32622 55074
rect 32674 55022 32676 55074
rect 32508 54404 32564 54414
rect 32508 54310 32564 54348
rect 32060 54238 32062 54290
rect 32114 54238 32116 54290
rect 32060 53732 32116 54238
rect 32620 53844 32676 55022
rect 32060 53666 32116 53676
rect 32508 53788 32676 53844
rect 33180 54514 33236 54526
rect 33180 54462 33182 54514
rect 33234 54462 33236 54514
rect 32060 53172 32116 53182
rect 31948 53170 32116 53172
rect 31948 53118 32062 53170
rect 32114 53118 32116 53170
rect 31948 53116 32116 53118
rect 32060 53106 32116 53116
rect 32284 53060 32340 53070
rect 30828 52946 30884 52958
rect 30828 52894 30830 52946
rect 30882 52894 30884 52946
rect 30828 52836 30884 52894
rect 30828 52770 30884 52780
rect 31948 52836 32004 52846
rect 31948 52742 32004 52780
rect 32284 52274 32340 53004
rect 32284 52222 32286 52274
rect 32338 52222 32340 52274
rect 32284 52210 32340 52222
rect 30548 51324 30660 51380
rect 32508 51380 32564 53788
rect 33068 53730 33124 53742
rect 33068 53678 33070 53730
rect 33122 53678 33124 53730
rect 32620 53620 32676 53630
rect 32620 53526 32676 53564
rect 33068 53620 33124 53678
rect 33068 53554 33124 53564
rect 33180 52948 33236 54462
rect 33404 54514 33460 54526
rect 33404 54462 33406 54514
rect 33458 54462 33460 54514
rect 33404 54404 33460 54462
rect 33404 54338 33460 54348
rect 33292 53844 33348 53854
rect 33292 53618 33348 53788
rect 33292 53566 33294 53618
rect 33346 53566 33348 53618
rect 33292 53554 33348 53566
rect 33404 52948 33460 52958
rect 33180 52854 33236 52892
rect 33292 52946 33460 52948
rect 33292 52894 33406 52946
rect 33458 52894 33460 52946
rect 33292 52892 33460 52894
rect 33292 52388 33348 52892
rect 33404 52882 33460 52892
rect 32844 52332 33348 52388
rect 32844 52276 32900 52332
rect 32844 52182 32900 52220
rect 30492 51314 30548 51324
rect 30380 51156 30436 51166
rect 30380 50596 30436 51100
rect 30380 50594 30548 50596
rect 30380 50542 30382 50594
rect 30434 50542 30548 50594
rect 30380 50540 30548 50542
rect 30380 50530 30436 50540
rect 30380 50036 30436 50046
rect 29260 49812 29316 49822
rect 29260 49698 29316 49756
rect 29260 49646 29262 49698
rect 29314 49646 29316 49698
rect 29260 49140 29316 49646
rect 29260 49074 29316 49084
rect 29596 49138 29652 49150
rect 29596 49086 29598 49138
rect 29650 49086 29652 49138
rect 29484 48356 29540 48366
rect 29036 48244 29092 48254
rect 29036 48150 29092 48188
rect 28588 48066 28644 48076
rect 29484 48020 29540 48300
rect 29484 47954 29540 47964
rect 29372 47458 29428 47470
rect 29372 47406 29374 47458
rect 29426 47406 29428 47458
rect 27916 46786 27972 46956
rect 27916 46734 27918 46786
rect 27970 46734 27972 46786
rect 27916 46722 27972 46734
rect 28140 47346 28196 47358
rect 28140 47294 28142 47346
rect 28194 47294 28196 47346
rect 27804 45950 27806 46002
rect 27858 45950 27860 46002
rect 27804 45938 27860 45950
rect 28140 45556 28196 47294
rect 29148 47346 29204 47358
rect 29148 47294 29150 47346
rect 29202 47294 29204 47346
rect 28812 46788 28868 46798
rect 28140 45490 28196 45500
rect 28252 46116 28308 46126
rect 27580 45278 27582 45330
rect 27634 45278 27636 45330
rect 27580 45266 27636 45278
rect 27468 44100 27524 44110
rect 27804 44100 27860 44110
rect 27524 44098 27860 44100
rect 27524 44046 27806 44098
rect 27858 44046 27860 44098
rect 27524 44044 27860 44046
rect 27468 44006 27524 44044
rect 27804 44034 27860 44044
rect 28252 43762 28308 46060
rect 28252 43710 28254 43762
rect 28306 43710 28308 43762
rect 28252 43698 28308 43710
rect 28364 45668 28420 45678
rect 28140 43540 28196 43550
rect 27468 43538 28196 43540
rect 27468 43486 28142 43538
rect 28194 43486 28196 43538
rect 27468 43484 28196 43486
rect 27020 42140 27300 42196
rect 27356 42642 27412 42654
rect 27356 42590 27358 42642
rect 27410 42590 27412 42642
rect 26908 41860 26964 41870
rect 26908 41186 26964 41804
rect 26908 41134 26910 41186
rect 26962 41134 26964 41186
rect 26908 41122 26964 41134
rect 27020 41188 27076 42140
rect 27356 42084 27412 42590
rect 27356 42018 27412 42028
rect 27244 41858 27300 41870
rect 27244 41806 27246 41858
rect 27298 41806 27300 41858
rect 27020 41122 27076 41132
rect 27132 41748 27188 41758
rect 27132 41186 27188 41692
rect 27132 41134 27134 41186
rect 27186 41134 27188 41186
rect 27132 40852 27188 41134
rect 27132 40786 27188 40796
rect 26684 40626 26852 40628
rect 26684 40574 26686 40626
rect 26738 40574 26852 40626
rect 26684 40572 26852 40574
rect 26684 40562 26740 40572
rect 27244 40516 27300 41806
rect 27356 40964 27412 40974
rect 27356 40628 27412 40908
rect 27356 40534 27412 40572
rect 27244 40450 27300 40460
rect 26460 39678 26462 39730
rect 26514 39678 26516 39730
rect 26460 39666 26516 39678
rect 26572 40404 26628 40414
rect 26012 38782 26014 38834
rect 26066 38782 26068 38834
rect 26012 38770 26068 38782
rect 26124 39620 26180 39630
rect 26124 38668 26180 39564
rect 26348 39284 26404 39294
rect 25788 38658 25844 38668
rect 25676 37538 25732 37548
rect 26012 38612 26180 38668
rect 26236 38724 26292 38762
rect 26236 38658 26292 38668
rect 26012 38052 26068 38612
rect 26236 38164 26292 38174
rect 26236 38070 26292 38108
rect 26012 37490 26068 37996
rect 26012 37438 26014 37490
rect 26066 37438 26068 37490
rect 26012 37426 26068 37438
rect 26124 38050 26180 38062
rect 26124 37998 26126 38050
rect 26178 37998 26180 38050
rect 25564 37326 25566 37378
rect 25618 37326 25620 37378
rect 25564 37156 25620 37326
rect 25564 37090 25620 37100
rect 25340 36642 25396 36652
rect 25788 37044 25844 37054
rect 25340 36484 25396 36494
rect 25340 36390 25396 36428
rect 25788 36482 25844 36988
rect 26124 36932 26180 37998
rect 26236 37380 26292 37390
rect 26236 37286 26292 37324
rect 26124 36866 26180 36876
rect 26012 36708 26068 36718
rect 26068 36652 26180 36708
rect 26012 36642 26068 36652
rect 25788 36430 25790 36482
rect 25842 36430 25844 36482
rect 25788 36418 25844 36430
rect 26012 36482 26068 36494
rect 26012 36430 26014 36482
rect 26066 36430 26068 36482
rect 25676 35924 25732 35934
rect 25732 35868 25844 35924
rect 25676 35858 25732 35868
rect 25228 35646 25230 35698
rect 25282 35646 25284 35698
rect 25228 35634 25284 35646
rect 25340 35812 25396 35822
rect 25340 35586 25396 35756
rect 25340 35534 25342 35586
rect 25394 35534 25396 35586
rect 25340 35522 25396 35534
rect 25452 35810 25508 35822
rect 25452 35758 25454 35810
rect 25506 35758 25508 35810
rect 25340 35252 25396 35262
rect 25228 34914 25284 34926
rect 25228 34862 25230 34914
rect 25282 34862 25284 34914
rect 25228 33460 25284 34862
rect 25340 34802 25396 35196
rect 25452 34916 25508 35758
rect 25452 34850 25508 34860
rect 25340 34750 25342 34802
rect 25394 34750 25396 34802
rect 25340 34738 25396 34750
rect 25228 33394 25284 33404
rect 25340 34130 25396 34142
rect 25340 34078 25342 34130
rect 25394 34078 25396 34130
rect 25340 33684 25396 34078
rect 25004 31950 25006 32002
rect 25058 31950 25060 32002
rect 25004 31938 25060 31950
rect 25116 33348 25172 33358
rect 25116 33236 25172 33292
rect 25228 33236 25284 33246
rect 25116 33234 25284 33236
rect 25116 33182 25230 33234
rect 25282 33182 25284 33234
rect 25116 33180 25284 33182
rect 25004 31780 25060 31790
rect 25116 31780 25172 33180
rect 25228 33170 25284 33180
rect 25340 33236 25396 33628
rect 25340 33170 25396 33180
rect 25564 34130 25620 34142
rect 25564 34078 25566 34130
rect 25618 34078 25620 34130
rect 25004 31778 25172 31780
rect 25004 31726 25006 31778
rect 25058 31726 25172 31778
rect 25004 31724 25172 31726
rect 25340 32564 25396 32574
rect 25004 31714 25060 31724
rect 25228 31668 25284 31678
rect 25116 31666 25284 31668
rect 25116 31614 25230 31666
rect 25282 31614 25284 31666
rect 25116 31612 25284 31614
rect 25116 30210 25172 31612
rect 25228 31602 25284 31612
rect 25340 30882 25396 32508
rect 25340 30830 25342 30882
rect 25394 30830 25396 30882
rect 25340 30818 25396 30830
rect 25564 32452 25620 34078
rect 25564 30660 25620 32396
rect 25452 30604 25620 30660
rect 25676 33346 25732 33358
rect 25676 33294 25678 33346
rect 25730 33294 25732 33346
rect 25676 30660 25732 33294
rect 25788 31220 25844 35868
rect 26012 35364 26068 36430
rect 26012 35298 26068 35308
rect 26124 34802 26180 36652
rect 26124 34750 26126 34802
rect 26178 34750 26180 34802
rect 26124 33906 26180 34750
rect 26236 35252 26292 35262
rect 26236 34244 26292 35196
rect 26348 35028 26404 39228
rect 26572 38948 26628 40348
rect 26684 39620 26740 39630
rect 26684 39284 26740 39564
rect 27020 39618 27076 39630
rect 27020 39566 27022 39618
rect 27074 39566 27076 39618
rect 27020 39396 27076 39566
rect 27132 39508 27188 39518
rect 27132 39414 27188 39452
rect 27020 39330 27076 39340
rect 26684 39218 26740 39228
rect 26684 38948 26740 38958
rect 26460 38946 26740 38948
rect 26460 38894 26686 38946
rect 26738 38894 26740 38946
rect 26460 38892 26740 38894
rect 26460 37044 26516 38892
rect 26684 38882 26740 38892
rect 27132 38948 27188 38958
rect 26908 38836 26964 38846
rect 26908 38742 26964 38780
rect 27132 38834 27188 38892
rect 27132 38782 27134 38834
rect 27186 38782 27188 38834
rect 27132 38770 27188 38782
rect 26572 38722 26628 38734
rect 26572 38670 26574 38722
rect 26626 38670 26628 38722
rect 26572 38276 26628 38670
rect 27468 38668 27524 43484
rect 28140 43474 28196 43484
rect 27804 42754 27860 42766
rect 27804 42702 27806 42754
rect 27858 42702 27860 42754
rect 27804 41748 27860 42702
rect 28252 42756 28308 42766
rect 28364 42756 28420 45612
rect 28700 45220 28756 45230
rect 28700 45126 28756 45164
rect 28476 44434 28532 44446
rect 28476 44382 28478 44434
rect 28530 44382 28532 44434
rect 28476 44212 28532 44382
rect 28476 44146 28532 44156
rect 28588 43538 28644 43550
rect 28588 43486 28590 43538
rect 28642 43486 28644 43538
rect 28588 43204 28644 43486
rect 28588 43138 28644 43148
rect 28364 42700 28532 42756
rect 27916 42644 27972 42654
rect 27916 42082 27972 42588
rect 27916 42030 27918 42082
rect 27970 42030 27972 42082
rect 27916 42018 27972 42030
rect 27804 41682 27860 41692
rect 28252 41410 28308 42700
rect 28364 42530 28420 42542
rect 28364 42478 28366 42530
rect 28418 42478 28420 42530
rect 28364 41748 28420 42478
rect 28364 41682 28420 41692
rect 28252 41358 28254 41410
rect 28306 41358 28308 41410
rect 28252 41346 28308 41358
rect 28476 41412 28532 42700
rect 28476 41356 28644 41412
rect 27916 41300 27972 41310
rect 27916 41206 27972 41244
rect 28364 41186 28420 41198
rect 28364 41134 28366 41186
rect 28418 41134 28420 41186
rect 27692 40852 27748 40862
rect 27580 40740 27636 40750
rect 27580 39730 27636 40684
rect 27692 40626 27748 40796
rect 27692 40574 27694 40626
rect 27746 40574 27748 40626
rect 27692 40562 27748 40574
rect 27580 39678 27582 39730
rect 27634 39678 27636 39730
rect 27580 39666 27636 39678
rect 27804 40516 27860 40526
rect 27804 39172 27860 40460
rect 28364 40404 28420 41134
rect 28364 40338 28420 40348
rect 28476 41188 28532 41198
rect 27916 40292 27972 40302
rect 27916 39842 27972 40236
rect 28252 40180 28308 40190
rect 27916 39790 27918 39842
rect 27970 39790 27972 39842
rect 27916 39778 27972 39790
rect 28028 39956 28084 39966
rect 28028 39842 28084 39900
rect 28028 39790 28030 39842
rect 28082 39790 28084 39842
rect 27580 39116 27860 39172
rect 27580 39058 27636 39116
rect 27580 39006 27582 39058
rect 27634 39006 27636 39058
rect 27580 38994 27636 39006
rect 27916 38948 27972 38958
rect 27916 38854 27972 38892
rect 27356 38612 27524 38668
rect 27692 38724 27748 38734
rect 28028 38668 28084 39790
rect 28252 39842 28308 40124
rect 28252 39790 28254 39842
rect 28306 39790 28308 39842
rect 28252 39620 28308 39790
rect 28252 39554 28308 39564
rect 28476 39618 28532 41132
rect 28588 40740 28644 41356
rect 28588 40402 28644 40684
rect 28588 40350 28590 40402
rect 28642 40350 28644 40402
rect 28588 40338 28644 40350
rect 28812 40402 28868 46732
rect 29148 43988 29204 47294
rect 29148 43922 29204 43932
rect 29260 46340 29316 46350
rect 29148 43652 29204 43662
rect 29148 43558 29204 43596
rect 28812 40350 28814 40402
rect 28866 40350 28868 40402
rect 28812 40338 28868 40350
rect 29148 41186 29204 41198
rect 29148 41134 29150 41186
rect 29202 41134 29204 41186
rect 29148 40964 29204 41134
rect 28476 39566 28478 39618
rect 28530 39566 28532 39618
rect 26572 38210 26628 38220
rect 27244 38388 27300 38398
rect 27244 37938 27300 38332
rect 27244 37886 27246 37938
rect 27298 37886 27300 37938
rect 27244 37874 27300 37886
rect 26796 37492 26852 37502
rect 26796 37398 26852 37436
rect 26572 37268 26628 37278
rect 26572 37174 26628 37212
rect 27244 37156 27300 37166
rect 27356 37156 27412 38612
rect 27692 37828 27748 38668
rect 27468 37268 27524 37278
rect 27524 37212 27636 37268
rect 27468 37202 27524 37212
rect 27020 37154 27412 37156
rect 27020 37102 27246 37154
rect 27298 37102 27412 37154
rect 27020 37100 27412 37102
rect 26460 36988 26852 37044
rect 26572 36820 26628 36830
rect 26460 35028 26516 35038
rect 26348 34972 26460 35028
rect 26460 34934 26516 34972
rect 26236 34130 26292 34188
rect 26236 34078 26238 34130
rect 26290 34078 26292 34130
rect 26236 34066 26292 34078
rect 26124 33854 26126 33906
rect 26178 33854 26180 33906
rect 26124 33842 26180 33854
rect 26460 33908 26516 33918
rect 26460 33234 26516 33852
rect 26572 33458 26628 36764
rect 26684 35586 26740 35598
rect 26684 35534 26686 35586
rect 26738 35534 26740 35586
rect 26684 35476 26740 35534
rect 26684 35410 26740 35420
rect 26796 35026 26852 36988
rect 26796 34974 26798 35026
rect 26850 34974 26852 35026
rect 26796 34962 26852 34974
rect 26908 36932 26964 36942
rect 26684 34916 26740 34926
rect 26684 34822 26740 34860
rect 26796 34132 26852 34142
rect 26572 33406 26574 33458
rect 26626 33406 26628 33458
rect 26572 33394 26628 33406
rect 26684 34076 26796 34132
rect 26460 33182 26462 33234
rect 26514 33182 26516 33234
rect 26460 33170 26516 33182
rect 26572 32676 26628 32686
rect 26124 31332 26180 31342
rect 25788 31218 26068 31220
rect 25788 31166 25790 31218
rect 25842 31166 26068 31218
rect 25788 31164 26068 31166
rect 25788 31154 25844 31164
rect 26012 30996 26068 31164
rect 26124 31218 26180 31276
rect 26124 31166 26126 31218
rect 26178 31166 26180 31218
rect 26124 31154 26180 31166
rect 26348 31220 26404 31230
rect 26348 31126 26404 31164
rect 26572 31218 26628 32620
rect 26572 31166 26574 31218
rect 26626 31166 26628 31218
rect 26572 31154 26628 31166
rect 26236 30996 26292 31006
rect 26012 30940 26180 30996
rect 25116 30158 25118 30210
rect 25170 30158 25172 30210
rect 25116 30100 25172 30158
rect 25228 30212 25284 30222
rect 25228 30118 25284 30156
rect 25116 30034 25172 30044
rect 25340 30098 25396 30110
rect 25340 30046 25342 30098
rect 25394 30046 25396 30098
rect 25340 29988 25396 30046
rect 25340 29922 25396 29932
rect 25116 28644 25172 28654
rect 25116 28550 25172 28588
rect 25452 28308 25508 30604
rect 25676 30594 25732 30604
rect 25900 30436 25956 30446
rect 25564 30210 25620 30222
rect 25564 30158 25566 30210
rect 25618 30158 25620 30210
rect 25564 29652 25620 30158
rect 25564 29586 25620 29596
rect 25900 29650 25956 30380
rect 26124 30436 26180 30940
rect 26236 30902 26292 30940
rect 26124 30380 26404 30436
rect 26012 29988 26068 29998
rect 26012 29894 26068 29932
rect 25900 29598 25902 29650
rect 25954 29598 25956 29650
rect 25900 29586 25956 29598
rect 25676 29316 25732 29326
rect 25452 28252 25620 28308
rect 25340 28084 25396 28094
rect 25340 27990 25396 28028
rect 24780 27246 24782 27298
rect 24834 27246 24836 27298
rect 24780 27234 24836 27246
rect 25228 27860 25284 27870
rect 24220 27188 24276 27198
rect 24220 27074 24276 27132
rect 24220 27022 24222 27074
rect 24274 27022 24276 27074
rect 24220 27010 24276 27022
rect 24444 27074 24500 27086
rect 24444 27022 24446 27074
rect 24498 27022 24500 27074
rect 24444 25844 24500 27022
rect 25228 27074 25284 27804
rect 25452 27858 25508 27870
rect 25452 27806 25454 27858
rect 25506 27806 25508 27858
rect 25452 27636 25508 27806
rect 25452 27570 25508 27580
rect 25228 27022 25230 27074
rect 25282 27022 25284 27074
rect 25228 27010 25284 27022
rect 25452 26292 25508 26302
rect 25452 26178 25508 26236
rect 25452 26126 25454 26178
rect 25506 26126 25508 26178
rect 25452 26114 25508 26126
rect 25564 26180 25620 28252
rect 25676 28082 25732 29260
rect 26012 29204 26068 29214
rect 26012 28644 26068 29148
rect 26012 28550 26068 28588
rect 25676 28030 25678 28082
rect 25730 28030 25732 28082
rect 25676 26964 25732 28030
rect 26124 27188 26180 30380
rect 26348 30322 26404 30380
rect 26348 30270 26350 30322
rect 26402 30270 26404 30322
rect 26348 30258 26404 30270
rect 26684 29988 26740 34076
rect 26796 34066 26852 34076
rect 26908 32452 26964 36876
rect 27020 36708 27076 37100
rect 27244 37090 27300 37100
rect 27468 37044 27524 37054
rect 27356 37042 27524 37044
rect 27356 36990 27470 37042
rect 27522 36990 27524 37042
rect 27356 36988 27524 36990
rect 27356 36932 27412 36988
rect 27468 36978 27524 36988
rect 27356 36866 27412 36876
rect 27580 36820 27636 37212
rect 27692 37266 27748 37772
rect 27692 37214 27694 37266
rect 27746 37214 27748 37266
rect 27692 37202 27748 37214
rect 27804 38612 28084 38668
rect 27468 36764 27636 36820
rect 27020 36652 27300 36708
rect 27132 35588 27188 35598
rect 27132 35364 27188 35532
rect 27132 35298 27188 35308
rect 27020 35140 27076 35150
rect 27020 34914 27076 35084
rect 27020 34862 27022 34914
rect 27074 34862 27076 34914
rect 27020 34132 27076 34862
rect 27132 35028 27188 35038
rect 27132 34914 27188 34972
rect 27132 34862 27134 34914
rect 27186 34862 27188 34914
rect 27132 34850 27188 34862
rect 27244 34692 27300 36652
rect 27468 35924 27524 36764
rect 27580 36596 27636 36606
rect 27580 36502 27636 36540
rect 27804 36036 27860 38612
rect 28364 38164 28420 38174
rect 28364 38070 28420 38108
rect 28252 37940 28308 37950
rect 28476 37940 28532 39566
rect 28700 39956 28756 39966
rect 28588 39172 28644 39182
rect 28588 38276 28644 39116
rect 28700 39058 28756 39900
rect 29148 39956 29204 40908
rect 29148 39890 29204 39900
rect 28700 39006 28702 39058
rect 28754 39006 28756 39058
rect 28700 38994 28756 39006
rect 29260 39620 29316 46284
rect 29372 46116 29428 47406
rect 29596 46900 29652 49086
rect 29820 48244 29876 48254
rect 29820 48150 29876 48188
rect 29596 46452 29652 46844
rect 30380 46564 30436 49980
rect 30492 48466 30548 50540
rect 30716 50370 30772 50382
rect 32396 50372 32452 50382
rect 30716 50318 30718 50370
rect 30770 50318 30772 50370
rect 30716 50036 30772 50318
rect 30716 49970 30772 49980
rect 32172 50316 32396 50372
rect 32172 49810 32228 50316
rect 32396 50278 32452 50316
rect 32172 49758 32174 49810
rect 32226 49758 32228 49810
rect 32172 49746 32228 49758
rect 30492 48414 30494 48466
rect 30546 48414 30548 48466
rect 30492 48402 30548 48414
rect 31388 49698 31444 49710
rect 31388 49646 31390 49698
rect 31442 49646 31444 49698
rect 31388 48466 31444 49646
rect 31836 49700 31892 49710
rect 31724 48914 31780 48926
rect 31724 48862 31726 48914
rect 31778 48862 31780 48914
rect 31724 48580 31780 48862
rect 31724 48514 31780 48524
rect 31388 48414 31390 48466
rect 31442 48414 31444 48466
rect 31388 48402 31444 48414
rect 30828 48354 30884 48366
rect 30828 48302 30830 48354
rect 30882 48302 30884 48354
rect 30828 48244 30884 48302
rect 31500 48356 31556 48366
rect 31500 48262 31556 48300
rect 31724 48356 31780 48366
rect 31836 48356 31892 49644
rect 32508 49252 32564 51324
rect 33516 52162 33572 55244
rect 33628 55206 33684 55244
rect 34300 55186 34356 55198
rect 34300 55134 34302 55186
rect 34354 55134 34356 55186
rect 33964 54740 34020 54750
rect 34300 54740 34356 55134
rect 33964 54738 34356 54740
rect 33964 54686 33966 54738
rect 34018 54686 34356 54738
rect 33964 54684 34356 54686
rect 33964 54674 34020 54684
rect 34748 54628 34804 54638
rect 34860 54628 34916 56142
rect 36764 56194 36820 56252
rect 39340 56306 39396 56590
rect 39340 56254 39342 56306
rect 39394 56254 39396 56306
rect 39340 56242 39396 56254
rect 40124 56642 40180 56654
rect 40124 56590 40126 56642
rect 40178 56590 40180 56642
rect 36764 56142 36766 56194
rect 36818 56142 36820 56194
rect 36764 56130 36820 56142
rect 37100 56194 37156 56206
rect 37100 56142 37102 56194
rect 37154 56142 37156 56194
rect 35196 55692 35460 55702
rect 35252 55636 35300 55692
rect 35356 55636 35404 55692
rect 35196 55626 35460 55636
rect 36428 55412 36484 55422
rect 36428 55410 36708 55412
rect 36428 55358 36430 55410
rect 36482 55358 36708 55410
rect 36428 55356 36708 55358
rect 36428 55346 36484 55356
rect 36428 54740 36484 54750
rect 34748 54626 34916 54628
rect 34748 54574 34750 54626
rect 34802 54574 34916 54626
rect 34748 54572 34916 54574
rect 36316 54738 36484 54740
rect 36316 54686 36430 54738
rect 36482 54686 36484 54738
rect 36316 54684 36484 54686
rect 36316 54628 36372 54684
rect 36428 54674 36484 54684
rect 34748 54562 34804 54572
rect 36316 54562 36372 54572
rect 36652 54626 36708 55356
rect 37100 55298 37156 56142
rect 39788 56194 39844 56206
rect 39788 56142 39790 56194
rect 39842 56142 39844 56194
rect 37100 55246 37102 55298
rect 37154 55246 37156 55298
rect 37100 55234 37156 55246
rect 37996 55970 38052 55982
rect 37996 55918 37998 55970
rect 38050 55918 38052 55970
rect 37324 55186 37380 55198
rect 37324 55134 37326 55186
rect 37378 55134 37380 55186
rect 36652 54574 36654 54626
rect 36706 54574 36708 54626
rect 33964 54514 34020 54526
rect 33964 54462 33966 54514
rect 34018 54462 34020 54514
rect 33964 54404 34020 54462
rect 33964 54338 34020 54348
rect 34412 54402 34468 54414
rect 34412 54350 34414 54402
rect 34466 54350 34468 54402
rect 33628 54290 33684 54302
rect 33628 54238 33630 54290
rect 33682 54238 33684 54290
rect 33628 53844 33684 54238
rect 33628 52946 33684 53788
rect 33964 53172 34020 53182
rect 34412 53172 34468 54350
rect 36316 54404 36372 54414
rect 36316 54310 36372 54348
rect 35196 54124 35460 54134
rect 35252 54068 35300 54124
rect 35356 54068 35404 54124
rect 35196 54058 35460 54068
rect 33964 53170 34244 53172
rect 33964 53118 33966 53170
rect 34018 53118 34244 53170
rect 33964 53116 34244 53118
rect 33964 53106 34020 53116
rect 33628 52894 33630 52946
rect 33682 52894 33684 52946
rect 33628 52882 33684 52894
rect 33964 52948 34020 52958
rect 33964 52854 34020 52892
rect 34188 52274 34244 53116
rect 34188 52222 34190 52274
rect 34242 52222 34244 52274
rect 34188 52210 34244 52222
rect 33516 52110 33518 52162
rect 33570 52110 33572 52162
rect 32396 49196 32564 49252
rect 32956 50372 33012 50382
rect 31724 48354 31892 48356
rect 31724 48302 31726 48354
rect 31778 48302 31892 48354
rect 31724 48300 31892 48302
rect 32172 48356 32228 48366
rect 31724 48290 31780 48300
rect 31164 48244 31220 48254
rect 30828 48242 31220 48244
rect 30828 48190 31166 48242
rect 31218 48190 31220 48242
rect 30828 48188 31220 48190
rect 30940 48020 30996 48030
rect 30940 47458 30996 47964
rect 30940 47406 30942 47458
rect 30994 47406 30996 47458
rect 30940 47394 30996 47406
rect 31164 47236 31220 48188
rect 32172 48130 32228 48300
rect 32172 48078 32174 48130
rect 32226 48078 32228 48130
rect 31500 47908 31556 47918
rect 31276 47460 31332 47470
rect 31276 47366 31332 47404
rect 31164 47170 31220 47180
rect 30380 46498 30436 46508
rect 31164 46676 31220 46686
rect 29596 46386 29652 46396
rect 29372 46050 29428 46060
rect 29372 45890 29428 45902
rect 29372 45838 29374 45890
rect 29426 45838 29428 45890
rect 29372 45332 29428 45838
rect 29372 45266 29428 45276
rect 29484 45778 29540 45790
rect 29484 45726 29486 45778
rect 29538 45726 29540 45778
rect 29372 44434 29428 44446
rect 29372 44382 29374 44434
rect 29426 44382 29428 44434
rect 29372 42756 29428 44382
rect 29372 42662 29428 42700
rect 29372 42196 29428 42206
rect 29484 42196 29540 45726
rect 29932 45108 29988 45118
rect 29932 45106 30212 45108
rect 29932 45054 29934 45106
rect 29986 45054 30212 45106
rect 29932 45052 30212 45054
rect 29932 45042 29988 45052
rect 30156 44548 30212 45052
rect 29596 44322 29652 44334
rect 29596 44270 29598 44322
rect 29650 44270 29652 44322
rect 29596 42308 29652 44270
rect 30044 44324 30100 44334
rect 29932 44210 29988 44222
rect 29932 44158 29934 44210
rect 29986 44158 29988 44210
rect 29932 43428 29988 44158
rect 29932 43362 29988 43372
rect 30044 42978 30100 44268
rect 30044 42926 30046 42978
rect 30098 42926 30100 42978
rect 30044 42914 30100 42926
rect 29932 42756 29988 42766
rect 29932 42754 30100 42756
rect 29932 42702 29934 42754
rect 29986 42702 30100 42754
rect 29932 42700 30100 42702
rect 29932 42690 29988 42700
rect 29596 42252 29988 42308
rect 29372 42194 29540 42196
rect 29372 42142 29374 42194
rect 29426 42142 29540 42194
rect 29372 42140 29540 42142
rect 29372 42130 29428 42140
rect 29596 41972 29652 41982
rect 29596 41878 29652 41916
rect 29932 41970 29988 42252
rect 29932 41918 29934 41970
rect 29986 41918 29988 41970
rect 29372 41186 29428 41198
rect 29372 41134 29374 41186
rect 29426 41134 29428 41186
rect 29372 40180 29428 41134
rect 29596 41188 29652 41198
rect 29596 41094 29652 41132
rect 29372 40114 29428 40124
rect 29484 40628 29540 40638
rect 29484 40292 29540 40572
rect 29484 39730 29540 40236
rect 29484 39678 29486 39730
rect 29538 39678 29540 39730
rect 29484 39666 29540 39678
rect 29260 39058 29316 39564
rect 29260 39006 29262 39058
rect 29314 39006 29316 39058
rect 29260 38994 29316 39006
rect 28588 38210 28644 38220
rect 28140 37938 28308 37940
rect 28140 37886 28254 37938
rect 28306 37886 28308 37938
rect 28140 37884 28308 37886
rect 27916 37156 27972 37166
rect 27916 37062 27972 37100
rect 27916 36932 27972 36942
rect 28140 36932 28196 37884
rect 28252 37874 28308 37884
rect 28364 37884 28532 37940
rect 28588 38050 28644 38062
rect 28588 37998 28590 38050
rect 28642 37998 28644 38050
rect 28364 37044 28420 37884
rect 27972 36876 28196 36932
rect 28252 36988 28420 37044
rect 28476 37154 28532 37166
rect 28476 37102 28478 37154
rect 28530 37102 28532 37154
rect 27916 36866 27972 36876
rect 28028 36372 28084 36382
rect 28028 36258 28084 36316
rect 28028 36206 28030 36258
rect 28082 36206 28084 36258
rect 28028 36148 28084 36206
rect 28252 36148 28308 36988
rect 28476 36484 28532 37102
rect 28588 37156 28644 37998
rect 29820 38050 29876 38062
rect 29820 37998 29822 38050
rect 29874 37998 29876 38050
rect 28588 37090 28644 37100
rect 28700 37940 28756 37950
rect 28532 36428 28644 36484
rect 28476 36390 28532 36428
rect 28364 36372 28420 36382
rect 28364 36278 28420 36316
rect 28476 36260 28532 36270
rect 28476 36166 28532 36204
rect 28252 36092 28420 36148
rect 28028 36082 28084 36092
rect 27020 34066 27076 34076
rect 27132 34636 27300 34692
rect 27356 35922 27524 35924
rect 27356 35870 27470 35922
rect 27522 35870 27524 35922
rect 27356 35868 27524 35870
rect 27020 33348 27076 33358
rect 27020 32676 27076 33292
rect 27020 32610 27076 32620
rect 26908 32396 27076 32452
rect 26796 32338 26852 32350
rect 26796 32286 26798 32338
rect 26850 32286 26852 32338
rect 26796 31778 26852 32286
rect 26796 31726 26798 31778
rect 26850 31726 26852 31778
rect 26796 30212 26852 31726
rect 26796 30146 26852 30156
rect 26684 29932 26852 29988
rect 26572 29316 26628 29326
rect 26572 29314 26740 29316
rect 26572 29262 26574 29314
rect 26626 29262 26740 29314
rect 26572 29260 26740 29262
rect 26572 29250 26628 29260
rect 26684 28868 26740 29260
rect 26684 28802 26740 28812
rect 26348 28756 26404 28766
rect 26348 27860 26404 28700
rect 26460 27860 26516 27870
rect 26348 27858 26516 27860
rect 26348 27806 26462 27858
rect 26514 27806 26516 27858
rect 26348 27804 26516 27806
rect 26460 27748 26516 27804
rect 26684 27860 26740 27870
rect 26684 27766 26740 27804
rect 26460 27682 26516 27692
rect 26572 27188 26628 27198
rect 26124 27186 26628 27188
rect 26124 27134 26574 27186
rect 26626 27134 26628 27186
rect 26124 27132 26628 27134
rect 26124 27076 26180 27132
rect 25900 27074 26180 27076
rect 25900 27022 26126 27074
rect 26178 27022 26180 27074
rect 25900 27020 26180 27022
rect 25788 26964 25844 26974
rect 25676 26962 25844 26964
rect 25676 26910 25790 26962
rect 25842 26910 25844 26962
rect 25676 26908 25844 26910
rect 25788 26898 25844 26908
rect 25900 26514 25956 27020
rect 26124 27010 26180 27020
rect 25900 26462 25902 26514
rect 25954 26462 25956 26514
rect 25900 26450 25956 26462
rect 26460 26514 26516 27132
rect 26572 27122 26628 27132
rect 26460 26462 26462 26514
rect 26514 26462 26516 26514
rect 26460 26450 26516 26462
rect 26796 26292 26852 29932
rect 26908 29204 26964 29214
rect 26908 28754 26964 29148
rect 26908 28702 26910 28754
rect 26962 28702 26964 28754
rect 26908 28690 26964 28702
rect 27020 28082 27076 32396
rect 27132 31890 27188 34636
rect 27244 34018 27300 34030
rect 27244 33966 27246 34018
rect 27298 33966 27300 34018
rect 27244 33684 27300 33966
rect 27244 33618 27300 33628
rect 27356 33348 27412 35868
rect 27468 35858 27524 35868
rect 27580 35980 27860 36036
rect 27580 35700 27636 35980
rect 28252 35924 28308 35934
rect 27356 33282 27412 33292
rect 27468 35644 27636 35700
rect 27692 35922 28308 35924
rect 27692 35870 28254 35922
rect 28306 35870 28308 35922
rect 27692 35868 28308 35870
rect 28364 35924 28420 36092
rect 28476 35924 28532 35934
rect 28364 35922 28532 35924
rect 28364 35870 28478 35922
rect 28530 35870 28532 35922
rect 28364 35868 28532 35870
rect 27468 32676 27524 35644
rect 27580 35476 27636 35486
rect 27580 34914 27636 35420
rect 27692 35026 27748 35868
rect 27804 35700 27860 35710
rect 27804 35606 27860 35644
rect 28140 35698 28196 35710
rect 28140 35646 28142 35698
rect 28194 35646 28196 35698
rect 27692 34974 27694 35026
rect 27746 34974 27748 35026
rect 27692 34962 27748 34974
rect 27804 35364 27860 35374
rect 27580 34862 27582 34914
rect 27634 34862 27636 34914
rect 27580 34850 27636 34862
rect 27804 34914 27860 35308
rect 27804 34862 27806 34914
rect 27858 34862 27860 34914
rect 27804 34850 27860 34862
rect 28028 34692 28084 34702
rect 28028 34598 28084 34636
rect 28140 34356 28196 35646
rect 28252 34580 28308 35868
rect 28476 35858 28532 35868
rect 28476 35476 28532 35486
rect 28252 34524 28420 34580
rect 28028 34300 28196 34356
rect 28252 34356 28308 34366
rect 28028 34244 28084 34300
rect 27916 34242 28084 34244
rect 27916 34190 28030 34242
rect 28082 34190 28084 34242
rect 27916 34188 28084 34190
rect 27580 33908 27636 33918
rect 27580 33814 27636 33852
rect 27804 33684 27860 33694
rect 27804 33346 27860 33628
rect 27916 33458 27972 34188
rect 28028 34178 28084 34188
rect 28252 34242 28308 34300
rect 28252 34190 28254 34242
rect 28306 34190 28308 34242
rect 28252 34178 28308 34190
rect 28140 34130 28196 34142
rect 28140 34078 28142 34130
rect 28194 34078 28196 34130
rect 28140 34020 28196 34078
rect 28364 34020 28420 34524
rect 28140 33964 28420 34020
rect 27916 33406 27918 33458
rect 27970 33406 27972 33458
rect 27916 33394 27972 33406
rect 27804 33294 27806 33346
rect 27858 33294 27860 33346
rect 27692 33124 27748 33134
rect 27692 33030 27748 33068
rect 27132 31838 27134 31890
rect 27186 31838 27188 31890
rect 27132 31826 27188 31838
rect 27356 32620 27524 32676
rect 27580 32788 27636 32798
rect 27132 30884 27188 30894
rect 27132 30790 27188 30828
rect 27244 30770 27300 30782
rect 27244 30718 27246 30770
rect 27298 30718 27300 30770
rect 27132 30324 27188 30334
rect 27244 30324 27300 30718
rect 27132 30322 27300 30324
rect 27132 30270 27134 30322
rect 27186 30270 27300 30322
rect 27132 30268 27300 30270
rect 27132 30258 27188 30268
rect 27132 29652 27188 29662
rect 27132 29558 27188 29596
rect 27356 29540 27412 32620
rect 27580 31218 27636 32732
rect 27692 32564 27748 32574
rect 27692 32470 27748 32508
rect 27804 32450 27860 33294
rect 28028 33348 28084 33358
rect 28028 32788 28084 33292
rect 28028 32722 28084 32732
rect 28252 33236 28308 33246
rect 28140 32564 28196 32574
rect 27804 32398 27806 32450
rect 27858 32398 27860 32450
rect 27804 32386 27860 32398
rect 28028 32562 28196 32564
rect 28028 32510 28142 32562
rect 28194 32510 28196 32562
rect 28028 32508 28196 32510
rect 28028 32004 28084 32508
rect 28140 32498 28196 32508
rect 27804 31948 28084 32004
rect 28252 32004 28308 33180
rect 28476 32788 28532 35420
rect 28588 35028 28644 36428
rect 28700 36482 28756 37884
rect 29708 37828 29764 37838
rect 29708 37734 29764 37772
rect 29372 37716 29428 37726
rect 29036 37380 29092 37390
rect 29036 37286 29092 37324
rect 28700 36430 28702 36482
rect 28754 36430 28756 36482
rect 28700 36418 28756 36430
rect 29036 37156 29092 37166
rect 29372 37156 29428 37660
rect 29596 37492 29652 37502
rect 29596 37398 29652 37436
rect 29708 37492 29764 37502
rect 29820 37492 29876 37998
rect 29708 37490 29876 37492
rect 29708 37438 29710 37490
rect 29762 37438 29876 37490
rect 29708 37436 29876 37438
rect 29708 37426 29764 37436
rect 29484 37380 29540 37390
rect 29484 37286 29540 37324
rect 29820 37268 29876 37278
rect 29596 37266 29876 37268
rect 29596 37214 29822 37266
rect 29874 37214 29876 37266
rect 29596 37212 29876 37214
rect 29596 37156 29652 37212
rect 29820 37202 29876 37212
rect 29372 37100 29652 37156
rect 28812 35700 28868 35710
rect 28812 35606 28868 35644
rect 28588 34962 28644 34972
rect 28700 34692 28756 34702
rect 28700 34598 28756 34636
rect 28812 34018 28868 34030
rect 28812 33966 28814 34018
rect 28866 33966 28868 34018
rect 28812 33348 28868 33966
rect 28812 33282 28868 33292
rect 28924 32788 28980 32798
rect 28476 32786 28980 32788
rect 28476 32734 28926 32786
rect 28978 32734 28980 32786
rect 28476 32732 28980 32734
rect 28364 32676 28420 32686
rect 28364 32582 28420 32620
rect 28476 32674 28532 32732
rect 28924 32722 28980 32732
rect 28476 32622 28478 32674
rect 28530 32622 28532 32674
rect 28476 32610 28532 32622
rect 28924 32564 28980 32574
rect 28252 31948 28644 32004
rect 27804 31666 27860 31948
rect 28252 31780 28308 31790
rect 28140 31778 28308 31780
rect 28140 31726 28254 31778
rect 28306 31726 28308 31778
rect 28140 31724 28308 31726
rect 28028 31668 28084 31678
rect 27804 31614 27806 31666
rect 27858 31614 27860 31666
rect 27804 31602 27860 31614
rect 27916 31666 28084 31668
rect 27916 31614 28030 31666
rect 28082 31614 28084 31666
rect 27916 31612 28084 31614
rect 27916 31444 27972 31612
rect 28028 31602 28084 31612
rect 27580 31166 27582 31218
rect 27634 31166 27636 31218
rect 27468 30884 27524 30894
rect 27580 30884 27636 31166
rect 27468 30882 27636 30884
rect 27468 30830 27470 30882
rect 27522 30830 27636 30882
rect 27468 30828 27636 30830
rect 27692 31388 27972 31444
rect 27468 30818 27524 30828
rect 27692 30548 27748 31388
rect 27804 31220 27860 31230
rect 27804 31126 27860 31164
rect 27916 31220 27972 31230
rect 28140 31220 28196 31724
rect 28252 31714 28308 31724
rect 27916 31218 28196 31220
rect 27916 31166 27918 31218
rect 27970 31166 28196 31218
rect 27916 31164 28196 31166
rect 27916 31154 27972 31164
rect 27692 30482 27748 30492
rect 28028 30994 28084 31006
rect 28028 30942 28030 30994
rect 28082 30942 28084 30994
rect 28028 30884 28084 30942
rect 28028 30324 28084 30828
rect 28028 30258 28084 30268
rect 28364 30436 28420 30446
rect 28364 30322 28420 30380
rect 28364 30270 28366 30322
rect 28418 30270 28420 30322
rect 28364 30258 28420 30270
rect 27580 30212 27636 30222
rect 27356 29484 27524 29540
rect 27244 29426 27300 29438
rect 27244 29374 27246 29426
rect 27298 29374 27300 29426
rect 27244 28868 27300 29374
rect 27244 28802 27300 28812
rect 27356 29316 27412 29326
rect 27356 28756 27412 29260
rect 27356 28662 27412 28700
rect 27020 28030 27022 28082
rect 27074 28030 27076 28082
rect 27020 28018 27076 28030
rect 27356 27972 27412 27982
rect 27356 27878 27412 27916
rect 27468 27412 27524 29484
rect 26796 26226 26852 26236
rect 27020 27356 27524 27412
rect 27580 27858 27636 30156
rect 27916 29988 27972 29998
rect 27692 29652 27748 29662
rect 27692 29558 27748 29596
rect 27916 29426 27972 29932
rect 27916 29374 27918 29426
rect 27970 29374 27972 29426
rect 27804 29316 27860 29326
rect 27804 29222 27860 29260
rect 27916 28868 27972 29374
rect 28364 29428 28420 29438
rect 28364 29334 28420 29372
rect 27580 27806 27582 27858
rect 27634 27806 27636 27858
rect 24444 25778 24500 25788
rect 25340 25620 25396 25630
rect 25340 25506 25396 25564
rect 25340 25454 25342 25506
rect 25394 25454 25396 25506
rect 25340 25442 25396 25454
rect 25564 25506 25620 26124
rect 25564 25454 25566 25506
rect 25618 25454 25620 25506
rect 25564 25442 25620 25454
rect 24444 25172 24500 25182
rect 24220 24834 24276 24846
rect 24220 24782 24222 24834
rect 24274 24782 24276 24834
rect 24220 24724 24276 24782
rect 24220 24658 24276 24668
rect 24444 24722 24500 25116
rect 25788 24948 25844 24958
rect 25452 24892 25788 24948
rect 24444 24670 24446 24722
rect 24498 24670 24500 24722
rect 24108 24546 24164 24556
rect 24332 24276 24388 24286
rect 24332 24050 24388 24220
rect 24332 23998 24334 24050
rect 24386 23998 24388 24050
rect 24332 23986 24388 23998
rect 24444 24052 24500 24670
rect 25004 24724 25060 24734
rect 25060 24668 25172 24724
rect 25004 24658 25060 24668
rect 25116 24052 25172 24668
rect 25228 24612 25284 24622
rect 25228 24518 25284 24556
rect 25228 24052 25284 24062
rect 25116 24050 25284 24052
rect 25116 23998 25230 24050
rect 25282 23998 25284 24050
rect 25116 23996 25284 23998
rect 24444 23986 24500 23996
rect 25228 23986 25284 23996
rect 24780 23940 24836 23950
rect 24780 23846 24836 23884
rect 25452 23940 25508 24892
rect 25788 24854 25844 24892
rect 26236 24948 26292 24958
rect 26236 24854 26292 24892
rect 25788 24052 25844 24062
rect 25788 23958 25844 23996
rect 23996 23426 24052 23436
rect 21644 23314 21700 23324
rect 22204 23286 22260 23324
rect 22988 23380 23044 23390
rect 22988 23286 23044 23324
rect 25452 23378 25508 23884
rect 25452 23326 25454 23378
rect 25506 23326 25508 23378
rect 25452 23314 25508 23326
rect 21364 23212 21476 23268
rect 21308 23174 21364 23212
rect 27020 23156 27076 27356
rect 27132 27188 27188 27198
rect 27580 27188 27636 27806
rect 27132 27186 27636 27188
rect 27132 27134 27134 27186
rect 27186 27134 27636 27186
rect 27132 27132 27636 27134
rect 27804 28812 27972 28868
rect 27132 27122 27188 27132
rect 27804 26628 27860 28812
rect 28252 28756 28308 28766
rect 28140 28530 28196 28542
rect 28140 28478 28142 28530
rect 28194 28478 28196 28530
rect 27804 26562 27860 26572
rect 27916 28420 27972 28430
rect 28140 28420 28196 28478
rect 28252 28530 28308 28700
rect 28476 28756 28532 28766
rect 28476 28642 28532 28700
rect 28476 28590 28478 28642
rect 28530 28590 28532 28642
rect 28476 28578 28532 28590
rect 28252 28478 28254 28530
rect 28306 28478 28308 28530
rect 28252 28466 28308 28478
rect 27916 28418 28196 28420
rect 27916 28366 27918 28418
rect 27970 28366 28196 28418
rect 27916 28364 28196 28366
rect 27916 27860 27972 28364
rect 27132 25620 27188 25630
rect 27132 25526 27188 25564
rect 27020 23090 27076 23100
rect 27804 25284 27860 25294
rect 19068 22930 19348 22932
rect 19068 22878 19070 22930
rect 19122 22878 19348 22930
rect 19068 22876 19348 22878
rect 19068 22866 19124 22876
rect 27804 22708 27860 25228
rect 27916 22932 27972 27804
rect 28140 27748 28196 27758
rect 28140 27654 28196 27692
rect 28588 27300 28644 31948
rect 28924 31218 28980 32508
rect 28924 31166 28926 31218
rect 28978 31166 28980 31218
rect 28924 31154 28980 31166
rect 28700 30994 28756 31006
rect 28700 30942 28702 30994
rect 28754 30942 28756 30994
rect 28700 30436 28756 30942
rect 28700 30370 28756 30380
rect 28812 30882 28868 30894
rect 28812 30830 28814 30882
rect 28866 30830 28868 30882
rect 28812 29652 28868 30830
rect 28812 29596 28980 29652
rect 28812 29426 28868 29438
rect 28812 29374 28814 29426
rect 28866 29374 28868 29426
rect 28700 28420 28756 28430
rect 28812 28420 28868 29374
rect 28924 29428 28980 29596
rect 28924 29362 28980 29372
rect 29036 29202 29092 37100
rect 29260 36260 29316 36270
rect 29260 36166 29316 36204
rect 29260 35586 29316 35598
rect 29260 35534 29262 35586
rect 29314 35534 29316 35586
rect 29260 35140 29316 35534
rect 29260 35074 29316 35084
rect 29372 35252 29428 35262
rect 29372 35026 29428 35196
rect 29372 34974 29374 35026
rect 29426 34974 29428 35026
rect 29260 34356 29316 34366
rect 29260 34262 29316 34300
rect 29260 33236 29316 33246
rect 29260 33142 29316 33180
rect 29148 33124 29204 33134
rect 29148 31890 29204 33068
rect 29148 31838 29150 31890
rect 29202 31838 29204 31890
rect 29148 31826 29204 31838
rect 29372 31220 29428 34974
rect 29484 32564 29540 32574
rect 29596 32564 29652 37100
rect 29932 36820 29988 41918
rect 30044 41410 30100 42700
rect 30156 41972 30212 44492
rect 30828 44324 30884 44334
rect 30828 44230 30884 44268
rect 30604 44210 30660 44222
rect 30604 44158 30606 44210
rect 30658 44158 30660 44210
rect 30604 43764 30660 44158
rect 30604 43698 30660 43708
rect 31052 43428 31108 43438
rect 30268 42754 30324 42766
rect 30268 42702 30270 42754
rect 30322 42702 30324 42754
rect 30268 42532 30324 42702
rect 31052 42754 31108 43372
rect 31052 42702 31054 42754
rect 31106 42702 31108 42754
rect 31052 42690 31108 42702
rect 30268 42084 30324 42476
rect 30828 42642 30884 42654
rect 30828 42590 30830 42642
rect 30882 42590 30884 42642
rect 30828 42196 30884 42590
rect 30828 42130 30884 42140
rect 30492 42084 30548 42094
rect 30268 42082 30548 42084
rect 30268 42030 30494 42082
rect 30546 42030 30548 42082
rect 30268 42028 30548 42030
rect 30492 42018 30548 42028
rect 30156 41906 30212 41916
rect 30044 41358 30046 41410
rect 30098 41358 30100 41410
rect 30044 41346 30100 41358
rect 31052 41076 31108 41086
rect 31052 40982 31108 41020
rect 30380 40964 30436 40974
rect 30044 40852 30100 40862
rect 30044 40180 30100 40796
rect 30156 40404 30212 40414
rect 30156 40310 30212 40348
rect 30380 40290 30436 40908
rect 30380 40238 30382 40290
rect 30434 40238 30436 40290
rect 30380 40226 30436 40238
rect 30828 40402 30884 40414
rect 30828 40350 30830 40402
rect 30882 40350 30884 40402
rect 30828 40292 30884 40350
rect 31164 40292 31220 46620
rect 31500 43652 31556 47852
rect 32060 47572 32116 47582
rect 32060 47478 32116 47516
rect 31948 47348 32004 47358
rect 31836 45892 31892 45902
rect 31836 45798 31892 45836
rect 31724 45778 31780 45790
rect 31724 45726 31726 45778
rect 31778 45726 31780 45778
rect 31724 44212 31780 45726
rect 31724 44146 31780 44156
rect 31724 43652 31780 43662
rect 31500 43650 31724 43652
rect 31500 43598 31502 43650
rect 31554 43598 31724 43650
rect 31500 43596 31724 43598
rect 31948 43652 32004 47292
rect 32060 46004 32116 46014
rect 32060 45910 32116 45948
rect 32172 44548 32228 48078
rect 32396 47068 32452 49196
rect 32956 49140 33012 50316
rect 33516 50372 33572 52110
rect 34412 50428 34468 53116
rect 34524 53620 34580 53630
rect 34524 50708 34580 53564
rect 36652 53058 36708 54574
rect 37100 55076 37156 55086
rect 36988 53732 37044 53742
rect 36652 53006 36654 53058
rect 36706 53006 36708 53058
rect 36652 52994 36708 53006
rect 36764 53060 36820 53070
rect 36764 52966 36820 53004
rect 36540 52946 36596 52958
rect 36540 52894 36542 52946
rect 36594 52894 36596 52946
rect 36540 52836 36596 52894
rect 36988 52946 37044 53676
rect 36988 52894 36990 52946
rect 37042 52894 37044 52946
rect 36988 52882 37044 52894
rect 36316 52780 36540 52836
rect 35196 52556 35460 52566
rect 35252 52500 35300 52556
rect 35356 52500 35404 52556
rect 35196 52490 35460 52500
rect 36316 52274 36372 52780
rect 36540 52770 36596 52780
rect 36316 52222 36318 52274
rect 36370 52222 36372 52274
rect 36316 52210 36372 52222
rect 37100 51938 37156 55020
rect 37100 51886 37102 51938
rect 37154 51886 37156 51938
rect 35196 50988 35460 50998
rect 35252 50932 35300 50988
rect 35356 50932 35404 50988
rect 35196 50922 35460 50932
rect 37100 50708 37156 51886
rect 34524 50706 35140 50708
rect 34524 50654 34526 50706
rect 34578 50654 35140 50706
rect 34524 50652 35140 50654
rect 34524 50642 34580 50652
rect 35084 50594 35140 50652
rect 35084 50542 35086 50594
rect 35138 50542 35140 50594
rect 35084 50530 35140 50542
rect 37100 50594 37156 50652
rect 37100 50542 37102 50594
rect 37154 50542 37156 50594
rect 33516 50306 33572 50316
rect 34300 50372 34468 50428
rect 34860 50372 34916 50382
rect 33068 50036 33124 50046
rect 33068 49942 33124 49980
rect 34076 50036 34132 50046
rect 33292 49812 33348 49822
rect 33292 49718 33348 49756
rect 33740 49810 33796 49822
rect 33740 49758 33742 49810
rect 33794 49758 33796 49810
rect 33180 49700 33236 49710
rect 33180 49606 33236 49644
rect 32508 49138 33012 49140
rect 32508 49086 32958 49138
rect 33010 49086 33012 49138
rect 32508 49084 33012 49086
rect 32508 49026 32564 49084
rect 32956 49074 33012 49084
rect 33516 49138 33572 49150
rect 33516 49086 33518 49138
rect 33570 49086 33572 49138
rect 32508 48974 32510 49026
rect 32562 48974 32564 49026
rect 32508 48962 32564 48974
rect 33516 48692 33572 49086
rect 33516 48626 33572 48636
rect 33068 48580 33124 48590
rect 32844 48132 32900 48142
rect 32844 47570 32900 48076
rect 32844 47518 32846 47570
rect 32898 47518 32900 47570
rect 32844 47460 32900 47518
rect 32844 47394 32900 47404
rect 32396 47012 32676 47068
rect 32620 46676 32676 47012
rect 33068 47012 33124 48524
rect 33628 48244 33684 48254
rect 33292 48242 33684 48244
rect 33292 48190 33630 48242
rect 33682 48190 33684 48242
rect 33292 48188 33684 48190
rect 33292 48130 33348 48188
rect 33628 48178 33684 48188
rect 33292 48078 33294 48130
rect 33346 48078 33348 48130
rect 33180 47460 33236 47470
rect 33180 47366 33236 47404
rect 33292 47124 33348 48078
rect 33740 47460 33796 49758
rect 33292 47058 33348 47068
rect 33516 47458 33796 47460
rect 33516 47406 33742 47458
rect 33794 47406 33796 47458
rect 33516 47404 33796 47406
rect 33516 47346 33572 47404
rect 33740 47394 33796 47404
rect 33964 49588 34020 49598
rect 33516 47294 33518 47346
rect 33570 47294 33572 47346
rect 33068 46956 33236 47012
rect 32620 46582 32676 46620
rect 32732 46900 32788 46910
rect 33180 46900 33236 46956
rect 33404 46900 33460 46910
rect 33180 46898 33460 46900
rect 33180 46846 33406 46898
rect 33458 46846 33460 46898
rect 33180 46844 33460 46846
rect 32508 46564 32564 46574
rect 32508 45332 32564 46508
rect 32732 45890 32788 46844
rect 33404 46834 33460 46844
rect 33068 46676 33124 46686
rect 32844 46674 33124 46676
rect 32844 46622 33070 46674
rect 33122 46622 33124 46674
rect 32844 46620 33124 46622
rect 32844 46002 32900 46620
rect 33068 46610 33124 46620
rect 33292 46676 33348 46686
rect 32844 45950 32846 46002
rect 32898 45950 32900 46002
rect 32844 45938 32900 45950
rect 32956 46452 33012 46462
rect 32732 45838 32734 45890
rect 32786 45838 32788 45890
rect 32732 45826 32788 45838
rect 32956 45890 33012 46396
rect 32956 45838 32958 45890
rect 33010 45838 33012 45890
rect 32956 45826 33012 45838
rect 33292 45668 33348 46620
rect 33404 45892 33460 45902
rect 33516 45892 33572 47294
rect 33628 47236 33684 47246
rect 33628 46786 33684 47180
rect 33628 46734 33630 46786
rect 33682 46734 33684 46786
rect 33628 46722 33684 46734
rect 33740 47012 33796 47022
rect 33404 45890 33572 45892
rect 33404 45838 33406 45890
rect 33458 45838 33572 45890
rect 33404 45836 33572 45838
rect 33404 45826 33460 45836
rect 33516 45780 33572 45836
rect 33516 45714 33572 45724
rect 33740 46002 33796 46956
rect 33964 46676 34020 49532
rect 34076 47236 34132 49980
rect 34300 49588 34356 50372
rect 34524 50370 34916 50372
rect 34524 50318 34862 50370
rect 34914 50318 34916 50370
rect 34524 50316 34916 50318
rect 34300 49522 34356 49532
rect 34412 49810 34468 49822
rect 34412 49758 34414 49810
rect 34466 49758 34468 49810
rect 34188 48692 34244 48702
rect 34188 47458 34244 48636
rect 34300 47572 34356 47582
rect 34412 47572 34468 49758
rect 34300 47570 34468 47572
rect 34300 47518 34302 47570
rect 34354 47518 34468 47570
rect 34300 47516 34468 47518
rect 34300 47506 34356 47516
rect 34188 47406 34190 47458
rect 34242 47406 34244 47458
rect 34188 47394 34244 47406
rect 34412 47236 34468 47246
rect 34076 47234 34468 47236
rect 34076 47182 34414 47234
rect 34466 47182 34468 47234
rect 34076 47180 34468 47182
rect 34076 46900 34132 47180
rect 34412 47170 34468 47180
rect 34076 46834 34132 46844
rect 34524 46788 34580 50316
rect 34860 50306 34916 50316
rect 37100 50372 37156 50542
rect 34748 49810 34804 49822
rect 34748 49758 34750 49810
rect 34802 49758 34804 49810
rect 34748 49588 34804 49758
rect 35084 49810 35140 49822
rect 35084 49758 35086 49810
rect 35138 49758 35140 49810
rect 34860 49700 34916 49710
rect 34860 49606 34916 49644
rect 34748 49522 34804 49532
rect 34972 47460 35028 47470
rect 34972 47366 35028 47404
rect 35084 47460 35140 49758
rect 35420 49698 35476 49710
rect 35420 49646 35422 49698
rect 35474 49646 35476 49698
rect 35420 49588 35476 49646
rect 35420 49522 35476 49532
rect 35644 49700 35700 49710
rect 35196 49420 35460 49430
rect 35252 49364 35300 49420
rect 35356 49364 35404 49420
rect 35196 49354 35460 49364
rect 35644 49138 35700 49644
rect 35644 49086 35646 49138
rect 35698 49086 35700 49138
rect 35644 49074 35700 49086
rect 36428 49026 36484 49038
rect 36428 48974 36430 49026
rect 36482 48974 36484 49026
rect 36428 48804 36484 48974
rect 36428 48738 36484 48748
rect 37100 48802 37156 50316
rect 37100 48750 37102 48802
rect 37154 48750 37156 48802
rect 37100 48692 37156 48750
rect 37100 48626 37156 48636
rect 37324 51492 37380 55134
rect 37772 55076 37828 55086
rect 37772 54982 37828 55020
rect 37884 54292 37940 54302
rect 37996 54292 38052 55918
rect 38892 55970 38948 55982
rect 38892 55918 38894 55970
rect 38946 55918 38948 55970
rect 38892 55860 38948 55918
rect 38892 55794 38948 55804
rect 39788 55468 39844 56142
rect 40124 56194 40180 56590
rect 41020 56308 41076 59200
rect 41468 56308 41524 56318
rect 41020 56306 41524 56308
rect 41020 56254 41470 56306
rect 41522 56254 41524 56306
rect 41020 56252 41524 56254
rect 41468 56242 41524 56252
rect 43260 56308 43316 59200
rect 43260 56242 43316 56252
rect 44604 56308 44660 56318
rect 44604 56214 44660 56252
rect 40124 56142 40126 56194
rect 40178 56142 40180 56194
rect 40124 56130 40180 56142
rect 40460 56082 40516 56094
rect 40460 56030 40462 56082
rect 40514 56030 40516 56082
rect 40460 55860 40516 56030
rect 40460 55794 40516 55804
rect 43708 56082 43764 56094
rect 43708 56030 43710 56082
rect 43762 56030 43764 56082
rect 39228 55412 39844 55468
rect 39228 55410 39284 55412
rect 39228 55358 39230 55410
rect 39282 55358 39284 55410
rect 39228 55346 39284 55358
rect 43148 55410 43204 55422
rect 43148 55358 43150 55410
rect 43202 55358 43204 55410
rect 40348 55298 40404 55310
rect 40348 55246 40350 55298
rect 40402 55246 40404 55298
rect 38220 55074 38276 55086
rect 38220 55022 38222 55074
rect 38274 55022 38276 55074
rect 38220 54628 38276 55022
rect 38220 54562 38276 54572
rect 38556 55074 38612 55086
rect 38556 55022 38558 55074
rect 38610 55022 38612 55074
rect 38556 54514 38612 55022
rect 39116 55074 39172 55086
rect 39116 55022 39118 55074
rect 39170 55022 39172 55074
rect 39116 54740 39172 55022
rect 39900 55076 39956 55086
rect 39900 54982 39956 55020
rect 40348 55076 40404 55246
rect 40348 55010 40404 55020
rect 41020 55186 41076 55198
rect 41020 55134 41022 55186
rect 41074 55134 41076 55186
rect 39116 54674 39172 54684
rect 40348 54740 40404 54750
rect 40348 54646 40404 54684
rect 40796 54740 40852 54750
rect 38892 54628 38948 54638
rect 38892 54534 38948 54572
rect 38556 54462 38558 54514
rect 38610 54462 38612 54514
rect 38220 54402 38276 54414
rect 38220 54350 38222 54402
rect 38274 54350 38276 54402
rect 38220 54292 38276 54350
rect 38556 54292 38612 54462
rect 37940 54236 38612 54292
rect 37772 53620 37828 53630
rect 37884 53620 37940 54236
rect 38332 53730 38388 54236
rect 39452 53956 39508 53966
rect 38332 53678 38334 53730
rect 38386 53678 38388 53730
rect 38332 53666 38388 53678
rect 39116 53844 39172 53854
rect 37772 53618 37940 53620
rect 37772 53566 37774 53618
rect 37826 53566 37940 53618
rect 37772 53564 37940 53566
rect 38444 53620 38500 53630
rect 38780 53620 38836 53630
rect 38500 53618 38836 53620
rect 38500 53566 38782 53618
rect 38834 53566 38836 53618
rect 38500 53564 38836 53566
rect 37772 53554 37828 53564
rect 38108 53506 38164 53518
rect 38108 53454 38110 53506
rect 38162 53454 38164 53506
rect 37772 52948 37828 52958
rect 37772 52854 37828 52892
rect 37996 52948 38052 52958
rect 38108 52948 38164 53454
rect 38444 53170 38500 53564
rect 38780 53554 38836 53564
rect 39116 53618 39172 53788
rect 39116 53566 39118 53618
rect 39170 53566 39172 53618
rect 39116 53554 39172 53566
rect 38444 53118 38446 53170
rect 38498 53118 38500 53170
rect 38444 53106 38500 53118
rect 37996 52946 38164 52948
rect 37996 52894 37998 52946
rect 38050 52894 38164 52946
rect 37996 52892 38164 52894
rect 37996 52882 38052 52892
rect 37660 52836 37716 52846
rect 37660 52742 37716 52780
rect 37436 52722 37492 52734
rect 37436 52670 37438 52722
rect 37490 52670 37492 52722
rect 37436 52164 37492 52670
rect 37436 52098 37492 52108
rect 38108 51716 38164 52892
rect 38668 52274 38724 52286
rect 38668 52222 38670 52274
rect 38722 52222 38724 52274
rect 38332 52164 38388 52174
rect 38332 52070 38388 52108
rect 38108 51650 38164 51660
rect 38668 51604 38724 52222
rect 39228 52052 39284 52062
rect 39228 51958 39284 51996
rect 38668 51538 38724 51548
rect 35196 47852 35460 47862
rect 35252 47796 35300 47852
rect 35356 47796 35404 47852
rect 35196 47786 35460 47796
rect 35756 47796 35812 47806
rect 35756 47570 35812 47740
rect 37324 47796 37380 51436
rect 38444 51380 38500 51390
rect 37884 51268 37940 51278
rect 37884 50706 37940 51212
rect 38444 51156 38500 51324
rect 38780 51380 38836 51390
rect 38780 51286 38836 51324
rect 39004 51378 39060 51390
rect 39004 51326 39006 51378
rect 39058 51326 39060 51378
rect 38892 51268 38948 51278
rect 38892 51174 38948 51212
rect 38444 51090 38500 51100
rect 39004 51156 39060 51326
rect 39004 51090 39060 51100
rect 39228 51156 39284 51166
rect 39228 51062 39284 51100
rect 37884 50654 37886 50706
rect 37938 50654 37940 50706
rect 37884 50642 37940 50654
rect 38892 48804 38948 48814
rect 38780 48802 39284 48804
rect 38780 48750 38894 48802
rect 38946 48750 39284 48802
rect 38780 48748 39284 48750
rect 38556 48692 38612 48702
rect 38556 48354 38612 48636
rect 38556 48302 38558 48354
rect 38610 48302 38612 48354
rect 38556 48290 38612 48302
rect 37324 47730 37380 47740
rect 38332 47796 38388 47806
rect 35756 47518 35758 47570
rect 35810 47518 35812 47570
rect 35308 47460 35364 47470
rect 35084 47458 35364 47460
rect 35084 47406 35310 47458
rect 35362 47406 35364 47458
rect 35084 47404 35364 47406
rect 34412 46732 34580 46788
rect 34748 47346 34804 47358
rect 34748 47294 34750 47346
rect 34802 47294 34804 47346
rect 33964 46620 34132 46676
rect 33740 45950 33742 46002
rect 33794 45950 33796 46002
rect 33404 45668 33460 45678
rect 33292 45612 33404 45668
rect 33404 45602 33460 45612
rect 32508 45330 33236 45332
rect 32508 45278 32510 45330
rect 32562 45278 33236 45330
rect 32508 45276 33236 45278
rect 32508 45266 32564 45276
rect 33180 45218 33236 45276
rect 33180 45166 33182 45218
rect 33234 45166 33236 45218
rect 33180 45154 33236 45166
rect 33404 45218 33460 45230
rect 33404 45166 33406 45218
rect 33458 45166 33460 45218
rect 32172 44482 32228 44492
rect 32732 44436 32788 44446
rect 32620 44380 32732 44436
rect 32620 44098 32676 44380
rect 32732 44370 32788 44380
rect 33292 44322 33348 44334
rect 33292 44270 33294 44322
rect 33346 44270 33348 44322
rect 32620 44046 32622 44098
rect 32674 44046 32676 44098
rect 32620 44034 32676 44046
rect 32956 44212 33012 44222
rect 32060 43652 32116 43662
rect 31948 43650 32116 43652
rect 31948 43598 32062 43650
rect 32114 43598 32116 43650
rect 31948 43596 32116 43598
rect 31500 43586 31556 43596
rect 31724 43558 31780 43596
rect 32060 41972 32116 43596
rect 32620 43652 32676 43662
rect 32620 43558 32676 43596
rect 32956 42642 33012 44156
rect 33292 44212 33348 44270
rect 33292 44146 33348 44156
rect 33404 43876 33460 45166
rect 33740 45108 33796 45950
rect 33852 45108 33908 45118
rect 33740 45106 33908 45108
rect 33740 45054 33854 45106
rect 33906 45054 33908 45106
rect 33740 45052 33908 45054
rect 33852 45042 33908 45052
rect 33516 44882 33572 44894
rect 33516 44830 33518 44882
rect 33570 44830 33572 44882
rect 33516 44324 33572 44830
rect 33516 44258 33572 44268
rect 33404 43820 33572 43876
rect 33068 43652 33124 43662
rect 33068 43558 33124 43596
rect 33404 43652 33460 43662
rect 33404 43558 33460 43596
rect 33516 43316 33572 43820
rect 33516 43250 33572 43260
rect 33964 43538 34020 43550
rect 33964 43486 33966 43538
rect 34018 43486 34020 43538
rect 33516 42756 33572 42766
rect 33516 42662 33572 42700
rect 32956 42590 32958 42642
rect 33010 42590 33012 42642
rect 32844 42532 32900 42542
rect 32844 42438 32900 42476
rect 32060 41906 32116 41916
rect 32844 42084 32900 42094
rect 31276 41186 31332 41198
rect 31276 41134 31278 41186
rect 31330 41134 31332 41186
rect 31276 40516 31332 41134
rect 32844 40964 32900 42028
rect 32956 41186 33012 42590
rect 33964 42420 34020 43486
rect 33964 42354 34020 42364
rect 33516 41972 33572 41982
rect 33516 41878 33572 41916
rect 34076 41860 34132 46620
rect 34188 45890 34244 45902
rect 34188 45838 34190 45890
rect 34242 45838 34244 45890
rect 34188 45780 34244 45838
rect 34188 45714 34244 45724
rect 34412 44546 34468 46732
rect 34524 46562 34580 46574
rect 34524 46510 34526 46562
rect 34578 46510 34580 46562
rect 34524 46228 34580 46510
rect 34580 46172 34692 46228
rect 34524 46162 34580 46172
rect 34636 45890 34692 46172
rect 34748 46002 34804 47294
rect 35084 47236 35140 47404
rect 35308 47394 35364 47404
rect 35756 47460 35812 47518
rect 37772 47684 37828 47694
rect 37772 47572 37828 47628
rect 37772 47570 38164 47572
rect 37772 47518 37774 47570
rect 37826 47518 38164 47570
rect 37772 47516 38164 47518
rect 37772 47506 37828 47516
rect 35756 47394 35812 47404
rect 38108 47460 38164 47516
rect 38108 47366 38164 47404
rect 35084 47170 35140 47180
rect 35196 47234 35252 47246
rect 35196 47182 35198 47234
rect 35250 47182 35252 47234
rect 34748 45950 34750 46002
rect 34802 45950 34804 46002
rect 34748 45938 34804 45950
rect 34860 46900 34916 46910
rect 34636 45838 34638 45890
rect 34690 45838 34692 45890
rect 34636 45826 34692 45838
rect 34860 45890 34916 46844
rect 35196 46788 35252 47182
rect 35196 46722 35252 46732
rect 36652 46788 36708 46798
rect 36652 46694 36708 46732
rect 37324 46674 37380 46686
rect 37324 46622 37326 46674
rect 37378 46622 37380 46674
rect 35196 46284 35460 46294
rect 35252 46228 35300 46284
rect 35356 46228 35404 46284
rect 35196 46218 35460 46228
rect 34860 45838 34862 45890
rect 34914 45838 34916 45890
rect 34860 45826 34916 45838
rect 34412 44494 34414 44546
rect 34466 44494 34468 44546
rect 34188 44324 34244 44334
rect 34188 44230 34244 44268
rect 34412 42980 34468 44494
rect 34412 42914 34468 42924
rect 34524 45668 34580 45678
rect 34524 42532 34580 45612
rect 36988 44996 37044 45006
rect 37324 44996 37380 46622
rect 36988 44994 37380 44996
rect 36988 44942 36990 44994
rect 37042 44942 37380 44994
rect 36988 44940 37380 44942
rect 37548 44996 37604 45006
rect 35196 44716 35460 44726
rect 35252 44660 35300 44716
rect 35356 44660 35404 44716
rect 35196 44650 35460 44660
rect 34748 44548 34804 44558
rect 34748 44322 34804 44492
rect 35420 44548 35476 44558
rect 35420 44434 35476 44492
rect 35420 44382 35422 44434
rect 35474 44382 35476 44434
rect 35420 44370 35476 44382
rect 34748 44270 34750 44322
rect 34802 44270 34804 44322
rect 34748 44258 34804 44270
rect 36316 44324 36372 44334
rect 34972 44210 35028 44222
rect 34972 44158 34974 44210
rect 35026 44158 35028 44210
rect 34636 44098 34692 44110
rect 34636 44046 34638 44098
rect 34690 44046 34692 44098
rect 34636 43650 34692 44046
rect 34636 43598 34638 43650
rect 34690 43598 34692 43650
rect 34636 43586 34692 43598
rect 34972 43652 35028 44158
rect 34636 42532 34692 42542
rect 34524 42530 34692 42532
rect 34524 42478 34638 42530
rect 34690 42478 34692 42530
rect 34524 42476 34692 42478
rect 34076 41766 34132 41804
rect 34524 42082 34580 42094
rect 34524 42030 34526 42082
rect 34578 42030 34580 42082
rect 34524 41972 34580 42030
rect 34636 42084 34692 42476
rect 34972 42084 35028 43596
rect 35196 43148 35460 43158
rect 35252 43092 35300 43148
rect 35356 43092 35404 43148
rect 35196 43082 35460 43092
rect 35308 42980 35364 42990
rect 34636 42018 34692 42028
rect 34748 42082 35028 42084
rect 34748 42030 34974 42082
rect 35026 42030 35028 42082
rect 34748 42028 35028 42030
rect 34300 41748 34356 41758
rect 34188 41746 34356 41748
rect 34188 41694 34302 41746
rect 34354 41694 34356 41746
rect 34188 41692 34356 41694
rect 32956 41134 32958 41186
rect 33010 41134 33012 41186
rect 32956 41122 33012 41134
rect 33516 41188 33572 41198
rect 33516 41094 33572 41132
rect 33068 40964 33124 40974
rect 32844 40908 33012 40964
rect 31276 40450 31332 40460
rect 31388 40402 31444 40414
rect 31388 40350 31390 40402
rect 31442 40350 31444 40402
rect 31164 40236 31332 40292
rect 30044 40124 30212 40180
rect 30044 39620 30100 39630
rect 30044 39526 30100 39564
rect 30044 38164 30100 38174
rect 30044 38070 30100 38108
rect 30044 37266 30100 37278
rect 30044 37214 30046 37266
rect 30098 37214 30100 37266
rect 30044 37156 30100 37214
rect 30044 37090 30100 37100
rect 29932 36754 29988 36764
rect 29708 36260 29764 36270
rect 29708 36166 29764 36204
rect 29820 35252 29876 35262
rect 29708 35028 29764 35038
rect 29708 34354 29764 34972
rect 29820 34914 29876 35196
rect 30156 34916 30212 40124
rect 30268 39844 30324 39854
rect 30268 39750 30324 39788
rect 30604 39618 30660 39630
rect 30604 39566 30606 39618
rect 30658 39566 30660 39618
rect 30604 38948 30660 39566
rect 30828 39618 30884 40236
rect 30828 39566 30830 39618
rect 30882 39566 30884 39618
rect 30828 39554 30884 39566
rect 31052 39396 31108 39406
rect 30940 38948 30996 38958
rect 30604 38946 30996 38948
rect 30604 38894 30942 38946
rect 30994 38894 30996 38946
rect 30604 38892 30996 38894
rect 30940 38882 30996 38892
rect 31052 38668 31108 39340
rect 30828 38612 31108 38668
rect 31164 38834 31220 38846
rect 31164 38782 31166 38834
rect 31218 38782 31220 38834
rect 30492 38052 30548 38062
rect 30492 37958 30548 37996
rect 30604 37940 30660 37950
rect 30604 37846 30660 37884
rect 30492 37044 30548 37054
rect 30492 36950 30548 36988
rect 29820 34862 29822 34914
rect 29874 34862 29876 34914
rect 29820 34850 29876 34862
rect 30044 34860 30212 34916
rect 30492 35026 30548 35038
rect 30492 34974 30494 35026
rect 30546 34974 30548 35026
rect 29708 34302 29710 34354
rect 29762 34302 29764 34354
rect 29708 34290 29764 34302
rect 30044 33572 30100 34860
rect 30380 34692 30436 34702
rect 30268 34020 30324 34030
rect 30268 33926 30324 33964
rect 30044 33516 30212 33572
rect 29540 32508 29652 32564
rect 29484 32498 29540 32508
rect 29372 30994 29428 31164
rect 29708 31556 29764 31566
rect 29708 31220 29764 31500
rect 29708 31154 29764 31164
rect 29372 30942 29374 30994
rect 29426 30942 29428 30994
rect 29372 30930 29428 30942
rect 29260 29988 29316 29998
rect 29260 29894 29316 29932
rect 29596 29538 29652 29550
rect 29596 29486 29598 29538
rect 29650 29486 29652 29538
rect 29484 29428 29540 29438
rect 29036 29150 29038 29202
rect 29090 29150 29092 29202
rect 29036 29138 29092 29150
rect 29148 29426 29540 29428
rect 29148 29374 29486 29426
rect 29538 29374 29540 29426
rect 29148 29372 29540 29374
rect 29148 28756 29204 29372
rect 29484 29362 29540 29372
rect 29148 28642 29204 28700
rect 29596 29316 29652 29486
rect 29148 28590 29150 28642
rect 29202 28590 29204 28642
rect 29148 28578 29204 28590
rect 29260 28642 29316 28654
rect 29260 28590 29262 28642
rect 29314 28590 29316 28642
rect 28756 28364 28868 28420
rect 29260 28420 29316 28590
rect 29596 28642 29652 29260
rect 29596 28590 29598 28642
rect 29650 28590 29652 28642
rect 29596 28578 29652 28590
rect 29708 29428 29764 29438
rect 29708 28642 29764 29372
rect 30156 28866 30212 33516
rect 30268 33346 30324 33358
rect 30268 33294 30270 33346
rect 30322 33294 30324 33346
rect 30268 29652 30324 33294
rect 30380 31890 30436 34636
rect 30380 31838 30382 31890
rect 30434 31838 30436 31890
rect 30380 31826 30436 31838
rect 30492 31780 30548 34974
rect 30716 34692 30772 34702
rect 30716 34354 30772 34636
rect 30716 34302 30718 34354
rect 30770 34302 30772 34354
rect 30716 33346 30772 34302
rect 30716 33294 30718 33346
rect 30770 33294 30772 33346
rect 30716 33282 30772 33294
rect 30492 31724 30772 31780
rect 30268 29586 30324 29596
rect 30492 30322 30548 30334
rect 30492 30270 30494 30322
rect 30546 30270 30548 30322
rect 30492 30100 30548 30270
rect 30492 29204 30548 30044
rect 30492 29138 30548 29148
rect 30156 28814 30158 28866
rect 30210 28814 30212 28866
rect 30156 28802 30212 28814
rect 29708 28590 29710 28642
rect 29762 28590 29764 28642
rect 29708 28578 29764 28590
rect 28700 28354 28756 28364
rect 29260 28354 29316 28364
rect 29708 28084 29764 28094
rect 29708 27990 29764 28028
rect 30604 28084 30660 28094
rect 30604 27990 30660 28028
rect 30044 27860 30100 27870
rect 30044 27766 30100 27804
rect 28588 27234 28644 27244
rect 29148 27746 29204 27758
rect 29148 27694 29150 27746
rect 29202 27694 29204 27746
rect 29148 27300 29204 27694
rect 29148 27234 29204 27244
rect 30716 26908 30772 31724
rect 30828 28196 30884 38612
rect 31164 38500 31220 38782
rect 31276 38668 31332 40236
rect 31388 39284 31444 40350
rect 32172 40404 32228 40414
rect 32172 39730 32228 40348
rect 32172 39678 32174 39730
rect 32226 39678 32228 39730
rect 32172 39666 32228 39678
rect 31388 39218 31444 39228
rect 31500 39618 31556 39630
rect 31500 39566 31502 39618
rect 31554 39566 31556 39618
rect 31500 38668 31556 39566
rect 31724 39620 31780 39630
rect 31724 39618 31892 39620
rect 31724 39566 31726 39618
rect 31778 39566 31892 39618
rect 31724 39564 31892 39566
rect 31724 39554 31780 39564
rect 31724 38834 31780 38846
rect 31724 38782 31726 38834
rect 31778 38782 31780 38834
rect 31276 38612 31444 38668
rect 31500 38612 31668 38668
rect 31164 38434 31220 38444
rect 31276 38164 31332 38174
rect 31052 38052 31108 38062
rect 31052 37266 31108 37996
rect 31052 37214 31054 37266
rect 31106 37214 31108 37266
rect 31052 37202 31108 37214
rect 31276 37266 31332 38108
rect 31276 37214 31278 37266
rect 31330 37214 31332 37266
rect 31276 37202 31332 37214
rect 30940 36036 30996 36046
rect 30996 35980 31108 36036
rect 30940 35970 30996 35980
rect 30940 35252 30996 35262
rect 30940 34914 30996 35196
rect 30940 34862 30942 34914
rect 30994 34862 30996 34914
rect 30940 34850 30996 34862
rect 30940 31556 30996 31566
rect 30940 30212 30996 31500
rect 30940 30118 30996 30156
rect 31052 30100 31108 35980
rect 31388 33572 31444 38612
rect 31500 37492 31556 37502
rect 31500 37266 31556 37436
rect 31500 37214 31502 37266
rect 31554 37214 31556 37266
rect 31500 37202 31556 37214
rect 31612 35140 31668 38612
rect 31724 37828 31780 38782
rect 31836 38050 31892 39564
rect 32844 39508 32900 39518
rect 32396 38946 32452 38958
rect 32396 38894 32398 38946
rect 32450 38894 32452 38946
rect 32396 38668 32452 38894
rect 32508 38836 32564 38846
rect 32844 38836 32900 39452
rect 32508 38834 32900 38836
rect 32508 38782 32510 38834
rect 32562 38782 32900 38834
rect 32508 38780 32900 38782
rect 32508 38770 32564 38780
rect 31836 37998 31838 38050
rect 31890 37998 31892 38050
rect 31836 37986 31892 37998
rect 32284 38612 32452 38668
rect 32060 37940 32116 37950
rect 32060 37846 32116 37884
rect 32172 37938 32228 37950
rect 32172 37886 32174 37938
rect 32226 37886 32228 37938
rect 31724 37762 31780 37772
rect 32172 37828 32228 37886
rect 32172 37762 32228 37772
rect 31724 37492 31780 37502
rect 31724 36594 31780 37436
rect 32060 37492 32116 37502
rect 32284 37492 32340 38612
rect 32116 37436 32340 37492
rect 32396 38500 32452 38510
rect 32060 37398 32116 37436
rect 32284 37268 32340 37278
rect 32396 37268 32452 38444
rect 32844 38162 32900 38780
rect 32844 38110 32846 38162
rect 32898 38110 32900 38162
rect 32844 38052 32900 38110
rect 32844 37986 32900 37996
rect 32284 37266 32396 37268
rect 32284 37214 32286 37266
rect 32338 37214 32396 37266
rect 32284 37212 32396 37214
rect 32284 37202 32340 37212
rect 32396 37174 32452 37212
rect 32732 37828 32788 37838
rect 31948 37156 32004 37166
rect 31948 37062 32004 37100
rect 31724 36542 31726 36594
rect 31778 36542 31780 36594
rect 31724 36530 31780 36542
rect 32732 36482 32788 37772
rect 32732 36430 32734 36482
rect 32786 36430 32788 36482
rect 32284 36258 32340 36270
rect 32284 36206 32286 36258
rect 32338 36206 32340 36258
rect 31612 35074 31668 35084
rect 31724 35700 31780 35710
rect 31724 34804 31780 35644
rect 32284 35700 32340 36206
rect 32284 35634 32340 35644
rect 31724 34738 31780 34748
rect 32396 34914 32452 34926
rect 32396 34862 32398 34914
rect 32450 34862 32452 34914
rect 31388 33506 31444 33516
rect 32172 33572 32228 33582
rect 32172 33478 32228 33516
rect 32396 33572 32452 34862
rect 32732 34914 32788 36430
rect 32732 34862 32734 34914
rect 32786 34862 32788 34914
rect 32732 34850 32788 34862
rect 32396 33506 32452 33516
rect 32620 34690 32676 34702
rect 32620 34638 32622 34690
rect 32674 34638 32676 34690
rect 32172 32788 32228 32798
rect 31500 30324 31556 30334
rect 31500 30230 31556 30268
rect 31948 30212 32004 30222
rect 31948 30118 32004 30156
rect 31052 30034 31108 30044
rect 30828 28130 30884 28140
rect 32172 26908 32228 32732
rect 32620 31668 32676 34638
rect 32956 33572 33012 40908
rect 33068 40870 33124 40908
rect 34076 40740 34132 40750
rect 34076 40626 34132 40684
rect 34076 40574 34078 40626
rect 34130 40574 34132 40626
rect 34076 40562 34132 40574
rect 33964 39620 34020 39630
rect 34188 39620 34244 41692
rect 34300 41682 34356 41692
rect 34524 40740 34580 41916
rect 34636 41748 34692 41758
rect 34636 41654 34692 41692
rect 34748 41188 34804 42028
rect 34972 42018 35028 42028
rect 35196 42084 35252 42094
rect 35196 41990 35252 42028
rect 35084 41860 35140 41870
rect 34972 41804 35084 41860
rect 34748 41186 34916 41188
rect 34748 41134 34750 41186
rect 34802 41134 34916 41186
rect 34748 41132 34916 41134
rect 34748 41122 34804 41132
rect 34524 40626 34580 40684
rect 34524 40574 34526 40626
rect 34578 40574 34580 40626
rect 34524 40562 34580 40574
rect 34636 40628 34692 40638
rect 34636 40290 34692 40572
rect 34860 40516 34916 41132
rect 34972 41074 35028 41804
rect 35084 41794 35140 41804
rect 35308 41748 35364 42924
rect 35420 42194 35476 42206
rect 35420 42142 35422 42194
rect 35474 42142 35476 42194
rect 35420 41972 35476 42142
rect 35420 41906 35476 41916
rect 35756 41972 35812 41982
rect 35756 41970 36036 41972
rect 35756 41918 35758 41970
rect 35810 41918 36036 41970
rect 35756 41916 36036 41918
rect 35756 41906 35812 41916
rect 35420 41748 35476 41758
rect 35756 41748 35812 41758
rect 35308 41746 35700 41748
rect 35308 41694 35422 41746
rect 35474 41694 35700 41746
rect 35308 41692 35700 41694
rect 35420 41682 35476 41692
rect 35196 41580 35460 41590
rect 35252 41524 35300 41580
rect 35356 41524 35404 41580
rect 35196 41514 35460 41524
rect 35308 41412 35364 41422
rect 35644 41412 35700 41692
rect 35364 41356 35476 41412
rect 35308 41318 35364 41356
rect 34972 41022 34974 41074
rect 35026 41022 35028 41074
rect 34972 41010 35028 41022
rect 35308 41186 35364 41198
rect 35308 41134 35310 41186
rect 35362 41134 35364 41186
rect 35196 40962 35252 40974
rect 35196 40910 35198 40962
rect 35250 40910 35252 40962
rect 34972 40516 35028 40526
rect 34860 40514 35028 40516
rect 34860 40462 34974 40514
rect 35026 40462 35028 40514
rect 34860 40460 35028 40462
rect 34972 40450 35028 40460
rect 34636 40238 34638 40290
rect 34690 40238 34692 40290
rect 34636 40226 34692 40238
rect 35196 40292 35252 40910
rect 35308 40628 35364 41134
rect 35308 40562 35364 40572
rect 35308 40404 35364 40414
rect 35308 40310 35364 40348
rect 35420 40402 35476 41356
rect 35644 41346 35700 41356
rect 35756 41188 35812 41692
rect 35980 41298 36036 41916
rect 36204 41858 36260 41870
rect 36204 41806 36206 41858
rect 36258 41806 36260 41858
rect 36204 41300 36260 41806
rect 35980 41246 35982 41298
rect 36034 41246 36036 41298
rect 35980 41234 36036 41246
rect 36092 41244 36260 41300
rect 35420 40350 35422 40402
rect 35474 40350 35476 40402
rect 35420 40338 35476 40350
rect 35532 41132 35812 41188
rect 35532 40402 35588 41132
rect 35868 41076 35924 41086
rect 35532 40350 35534 40402
rect 35586 40350 35588 40402
rect 35532 40338 35588 40350
rect 35644 41074 35924 41076
rect 35644 41022 35870 41074
rect 35922 41022 35924 41074
rect 35644 41020 35924 41022
rect 35196 40226 35252 40236
rect 33964 39618 34244 39620
rect 33964 39566 33966 39618
rect 34018 39566 34244 39618
rect 33964 39564 34244 39566
rect 34300 40178 34356 40190
rect 34300 40126 34302 40178
rect 34354 40126 34356 40178
rect 34300 39618 34356 40126
rect 35532 40180 35588 40190
rect 35196 40012 35460 40022
rect 35252 39956 35300 40012
rect 35356 39956 35404 40012
rect 35196 39946 35460 39956
rect 34300 39566 34302 39618
rect 34354 39566 34356 39618
rect 33964 39554 34020 39564
rect 33740 39508 33796 39518
rect 33740 39414 33796 39452
rect 33628 39284 33684 39294
rect 33628 38722 33684 39228
rect 33628 38670 33630 38722
rect 33682 38670 33684 38722
rect 33628 38658 33684 38670
rect 34076 38668 34132 39564
rect 34300 38834 34356 39566
rect 34636 39508 34692 39518
rect 34412 39506 34692 39508
rect 34412 39454 34638 39506
rect 34690 39454 34692 39506
rect 34412 39452 34692 39454
rect 34412 38948 34468 39452
rect 34636 39442 34692 39452
rect 35308 38948 35364 38958
rect 35532 38948 35588 40124
rect 34412 38946 34580 38948
rect 34412 38894 34414 38946
rect 34466 38894 34580 38946
rect 34412 38892 34580 38894
rect 34412 38882 34468 38892
rect 34300 38782 34302 38834
rect 34354 38782 34356 38834
rect 34300 38724 34356 38782
rect 34076 38612 34244 38668
rect 34300 38658 34356 38668
rect 34188 38164 34244 38612
rect 34188 38070 34244 38108
rect 33292 38050 33348 38062
rect 33292 37998 33294 38050
rect 33346 37998 33348 38050
rect 33292 37940 33348 37998
rect 33180 36484 33236 36494
rect 33068 36428 33180 36484
rect 33068 34130 33124 36428
rect 33180 36390 33236 36428
rect 33180 35140 33236 35150
rect 33180 34802 33236 35084
rect 33180 34750 33182 34802
rect 33234 34750 33236 34802
rect 33180 34738 33236 34750
rect 33068 34078 33070 34130
rect 33122 34078 33124 34130
rect 33068 34066 33124 34078
rect 32620 31602 32676 31612
rect 32844 33516 33012 33572
rect 33292 33572 33348 37884
rect 33740 37828 33796 37838
rect 33740 37734 33796 37772
rect 34188 37268 34244 37278
rect 33964 37212 34188 37268
rect 33852 36260 33908 36270
rect 33852 36166 33908 36204
rect 33404 35922 33460 35934
rect 33404 35870 33406 35922
rect 33458 35870 33460 35922
rect 33404 35252 33460 35870
rect 33852 35812 33908 35822
rect 33964 35812 34020 37212
rect 34188 37174 34244 37212
rect 34412 36482 34468 36494
rect 34412 36430 34414 36482
rect 34466 36430 34468 36482
rect 34412 35924 34468 36430
rect 34412 35858 34468 35868
rect 33852 35810 34020 35812
rect 33852 35758 33854 35810
rect 33906 35758 34020 35810
rect 33852 35756 34020 35758
rect 33852 35746 33908 35756
rect 33404 35186 33460 35196
rect 34524 34916 34580 38892
rect 35308 38946 35588 38948
rect 35308 38894 35310 38946
rect 35362 38894 35588 38946
rect 35308 38892 35588 38894
rect 35308 38882 35364 38892
rect 34412 34860 34580 34916
rect 34636 38724 34692 38734
rect 32844 29988 32900 33516
rect 33292 33506 33348 33516
rect 34188 34018 34244 34030
rect 34188 33966 34190 34018
rect 34242 33966 34244 34018
rect 33180 33460 33236 33470
rect 32956 33236 33012 33246
rect 33180 33236 33236 33404
rect 32956 33234 33236 33236
rect 32956 33182 32958 33234
rect 33010 33182 33236 33234
rect 32956 33180 33236 33182
rect 32956 33170 33012 33180
rect 33180 32674 33236 33180
rect 33180 32622 33182 32674
rect 33234 32622 33236 32674
rect 33180 31666 33236 32622
rect 33404 33346 33460 33358
rect 33404 33294 33406 33346
rect 33458 33294 33460 33346
rect 33404 32676 33460 33294
rect 33852 33236 33908 33274
rect 33852 33170 33908 33180
rect 33404 32610 33460 32620
rect 33852 33012 33908 33022
rect 33852 31890 33908 32956
rect 33852 31838 33854 31890
rect 33906 31838 33908 31890
rect 33852 31826 33908 31838
rect 34076 32786 34132 32798
rect 34076 32734 34078 32786
rect 34130 32734 34132 32786
rect 33180 31614 33182 31666
rect 33234 31614 33236 31666
rect 33180 31602 33236 31614
rect 33740 31778 33796 31790
rect 33740 31726 33742 31778
rect 33794 31726 33796 31778
rect 33180 31220 33236 31230
rect 33180 31126 33236 31164
rect 33740 30996 33796 31726
rect 33740 30930 33796 30940
rect 32844 29922 32900 29932
rect 34076 26908 34132 32734
rect 34188 32564 34244 33966
rect 34188 31778 34244 32508
rect 34188 31726 34190 31778
rect 34242 31726 34244 31778
rect 34188 31714 34244 31726
rect 34300 33572 34356 33582
rect 34188 31108 34244 31118
rect 34188 29540 34244 31052
rect 34300 31106 34356 33516
rect 34300 31054 34302 31106
rect 34354 31054 34356 31106
rect 34300 30884 34356 31054
rect 34412 31108 34468 34860
rect 34636 34804 34692 38668
rect 35084 38724 35140 38734
rect 34748 37266 34804 37278
rect 34748 37214 34750 37266
rect 34802 37214 34804 37266
rect 34748 35476 34804 37214
rect 35084 37266 35140 38668
rect 35196 38444 35460 38454
rect 35252 38388 35300 38444
rect 35356 38388 35404 38444
rect 35196 38378 35460 38388
rect 35084 37214 35086 37266
rect 35138 37214 35140 37266
rect 35084 37202 35140 37214
rect 35196 36876 35460 36886
rect 35252 36820 35300 36876
rect 35356 36820 35404 36876
rect 35196 36810 35460 36820
rect 35532 35924 35588 38892
rect 35644 37268 35700 41020
rect 35868 41010 35924 41020
rect 36092 40962 36148 41244
rect 36092 40910 36094 40962
rect 36146 40910 36148 40962
rect 36092 40740 36148 40910
rect 36092 40674 36148 40684
rect 35756 40626 35812 40638
rect 35756 40574 35758 40626
rect 35810 40574 35812 40626
rect 35756 38948 35812 40574
rect 36316 40626 36372 44268
rect 36988 43540 37044 44940
rect 37548 44434 37604 44940
rect 38332 44884 38388 47740
rect 38444 47234 38500 47246
rect 38444 47182 38446 47234
rect 38498 47182 38500 47234
rect 38444 46788 38500 47182
rect 38780 47236 38836 48748
rect 38892 48738 38948 48748
rect 39228 48466 39284 48748
rect 39228 48414 39230 48466
rect 39282 48414 39284 48466
rect 39228 48402 39284 48414
rect 39452 48244 39508 53900
rect 40236 52162 40292 52174
rect 40236 52110 40238 52162
rect 40290 52110 40292 52162
rect 40012 51604 40068 51614
rect 40012 51510 40068 51548
rect 40236 51492 40292 52110
rect 40124 51490 40292 51492
rect 40124 51438 40238 51490
rect 40290 51438 40292 51490
rect 40124 51436 40292 51438
rect 39564 51378 39620 51390
rect 39564 51326 39566 51378
rect 39618 51326 39620 51378
rect 39564 51268 39620 51326
rect 39900 51268 39956 51278
rect 39564 51266 39956 51268
rect 39564 51214 39902 51266
rect 39954 51214 39956 51266
rect 39564 51212 39956 51214
rect 39900 51202 39956 51212
rect 40012 50708 40068 50718
rect 40124 50708 40180 51436
rect 40236 51426 40292 51436
rect 40012 50706 40180 50708
rect 40012 50654 40014 50706
rect 40066 50654 40180 50706
rect 40012 50652 40180 50654
rect 40348 51044 40404 51054
rect 40012 50642 40068 50652
rect 40012 48692 40068 48702
rect 39452 48178 39508 48188
rect 39564 48354 39620 48366
rect 39564 48302 39566 48354
rect 39618 48302 39620 48354
rect 38780 47170 38836 47180
rect 38892 47460 38948 47470
rect 38444 46722 38500 46732
rect 38668 47012 38724 47022
rect 38556 45892 38612 45902
rect 38556 45798 38612 45836
rect 38668 45890 38724 46956
rect 38892 46898 38948 47404
rect 39004 47460 39060 47470
rect 39004 47458 39396 47460
rect 39004 47406 39006 47458
rect 39058 47406 39396 47458
rect 39004 47404 39396 47406
rect 39004 47394 39060 47404
rect 38892 46846 38894 46898
rect 38946 46846 38948 46898
rect 38892 46564 38948 46846
rect 39116 47234 39172 47246
rect 39116 47182 39118 47234
rect 39170 47182 39172 47234
rect 39116 46900 39172 47182
rect 39228 47234 39284 47246
rect 39228 47182 39230 47234
rect 39282 47182 39284 47234
rect 39228 47012 39284 47182
rect 39228 46946 39284 46956
rect 39116 46834 39172 46844
rect 39340 46788 39396 47404
rect 39564 47348 39620 48302
rect 39452 47292 39620 47348
rect 39900 47570 39956 47582
rect 39900 47518 39902 47570
rect 39954 47518 39956 47570
rect 39452 47234 39508 47292
rect 39452 47182 39454 47234
rect 39506 47182 39508 47234
rect 39452 47012 39508 47182
rect 39788 47012 39844 47022
rect 39900 47012 39956 47518
rect 39452 46956 39732 47012
rect 39452 46788 39508 46798
rect 39340 46786 39508 46788
rect 39340 46734 39454 46786
rect 39506 46734 39508 46786
rect 39340 46732 39508 46734
rect 39116 46674 39172 46686
rect 39116 46622 39118 46674
rect 39170 46622 39172 46674
rect 39116 46564 39172 46622
rect 38892 46508 39172 46564
rect 38668 45838 38670 45890
rect 38722 45838 38724 45890
rect 38668 45826 38724 45838
rect 39452 45108 39508 46732
rect 39452 45042 39508 45052
rect 39564 46788 39620 46798
rect 38332 44828 38612 44884
rect 37548 44382 37550 44434
rect 37602 44382 37604 44434
rect 37548 44370 37604 44382
rect 38556 44434 38612 44828
rect 38556 44382 38558 44434
rect 38610 44382 38612 44434
rect 38556 44324 38612 44382
rect 38556 44258 38612 44268
rect 39004 44322 39060 44334
rect 39004 44270 39006 44322
rect 39058 44270 39060 44322
rect 37436 44212 37492 44222
rect 37436 44118 37492 44156
rect 36764 43428 36820 43438
rect 36652 43426 36820 43428
rect 36652 43374 36766 43426
rect 36818 43374 36820 43426
rect 36652 43372 36820 43374
rect 36316 40574 36318 40626
rect 36370 40574 36372 40626
rect 36316 40404 36372 40574
rect 36316 40338 36372 40348
rect 36428 43316 36484 43326
rect 35756 38882 35812 38892
rect 35868 40292 35924 40302
rect 35868 37378 35924 40236
rect 36428 40180 36484 43260
rect 36428 40114 36484 40124
rect 36652 38668 36708 43372
rect 36764 43362 36820 43372
rect 36988 42420 37044 43484
rect 37212 43428 37268 43438
rect 37212 43334 37268 43372
rect 38668 43428 38724 43438
rect 38668 42868 38724 43372
rect 39004 42868 39060 44270
rect 39116 44324 39172 44334
rect 39116 44230 39172 44268
rect 39564 44322 39620 46732
rect 39564 44270 39566 44322
rect 39618 44270 39620 44322
rect 39340 44098 39396 44110
rect 39340 44046 39342 44098
rect 39394 44046 39396 44098
rect 39340 43650 39396 44046
rect 39340 43598 39342 43650
rect 39394 43598 39396 43650
rect 39340 43586 39396 43598
rect 39452 43652 39508 43662
rect 39116 42868 39172 42878
rect 39004 42866 39172 42868
rect 39004 42814 39118 42866
rect 39170 42814 39172 42866
rect 39004 42812 39172 42814
rect 38668 42774 38724 42812
rect 39116 42802 39172 42812
rect 39228 42868 39284 42878
rect 38556 42756 38612 42766
rect 38556 42662 38612 42700
rect 39228 42754 39284 42812
rect 39228 42702 39230 42754
rect 39282 42702 39284 42754
rect 39228 42690 39284 42702
rect 39004 42644 39060 42654
rect 39004 42550 39060 42588
rect 39452 42642 39508 43596
rect 39564 43204 39620 44270
rect 39676 45106 39732 46956
rect 39844 46956 39956 47012
rect 40012 47460 40068 48636
rect 39788 46946 39844 46956
rect 40012 46898 40068 47404
rect 40012 46846 40014 46898
rect 40066 46846 40068 46898
rect 40012 46834 40068 46846
rect 40348 47012 40404 50988
rect 40460 50708 40516 50718
rect 40460 50614 40516 50652
rect 40348 46898 40404 46956
rect 40348 46846 40350 46898
rect 40402 46846 40404 46898
rect 40348 46834 40404 46846
rect 40796 46004 40852 54684
rect 40908 54740 40964 54750
rect 41020 54740 41076 55134
rect 40908 54738 41076 54740
rect 40908 54686 40910 54738
rect 40962 54686 41076 54738
rect 40908 54684 41076 54686
rect 41356 54740 41412 54750
rect 40908 54674 40964 54684
rect 41244 54628 41300 54638
rect 41132 54572 41244 54628
rect 40908 54516 40964 54526
rect 40908 53954 40964 54460
rect 40908 53902 40910 53954
rect 40962 53902 40964 53954
rect 40908 53890 40964 53902
rect 41020 54514 41076 54526
rect 41020 54462 41022 54514
rect 41074 54462 41076 54514
rect 41020 53842 41076 54462
rect 41020 53790 41022 53842
rect 41074 53790 41076 53842
rect 41020 53778 41076 53790
rect 41020 53172 41076 53182
rect 41020 52722 41076 53116
rect 41020 52670 41022 52722
rect 41074 52670 41076 52722
rect 41020 52658 41076 52670
rect 41132 52052 41188 54572
rect 41244 54562 41300 54572
rect 41356 54514 41412 54684
rect 41692 54628 41748 54638
rect 41692 54534 41748 54572
rect 41356 54462 41358 54514
rect 41410 54462 41412 54514
rect 41356 54450 41412 54462
rect 41244 54292 41300 54302
rect 41244 54290 41748 54292
rect 41244 54238 41246 54290
rect 41298 54238 41748 54290
rect 41244 54236 41748 54238
rect 41244 54226 41300 54236
rect 41692 53844 41748 54236
rect 42140 53844 42196 53854
rect 41244 53732 41300 53742
rect 41244 53638 41300 53676
rect 41580 53060 41636 53070
rect 41468 52948 41524 52958
rect 41356 52892 41468 52948
rect 41244 52052 41300 52062
rect 41020 52050 41300 52052
rect 41020 51998 41246 52050
rect 41298 51998 41300 52050
rect 41020 51996 41300 51998
rect 41020 51490 41076 51996
rect 41244 51986 41300 51996
rect 41356 52050 41412 52892
rect 41468 52882 41524 52892
rect 41580 52834 41636 53004
rect 41580 52782 41582 52834
rect 41634 52782 41636 52834
rect 41468 52722 41524 52734
rect 41468 52670 41470 52722
rect 41522 52670 41524 52722
rect 41468 52162 41524 52670
rect 41468 52110 41470 52162
rect 41522 52110 41524 52162
rect 41468 52098 41524 52110
rect 41356 51998 41358 52050
rect 41410 51998 41412 52050
rect 41356 51986 41412 51998
rect 41580 51828 41636 52782
rect 41468 51772 41636 51828
rect 41692 52386 41748 53788
rect 42028 53842 42196 53844
rect 42028 53790 42142 53842
rect 42194 53790 42196 53842
rect 42028 53788 42196 53790
rect 41916 53060 41972 53070
rect 41916 52946 41972 53004
rect 41916 52894 41918 52946
rect 41970 52894 41972 52946
rect 41916 52882 41972 52894
rect 42028 52724 42084 53788
rect 42140 53778 42196 53788
rect 43148 53732 43204 55358
rect 43596 55076 43652 55086
rect 43708 55076 43764 56030
rect 45500 55412 45556 59200
rect 47740 56308 47796 59200
rect 47740 56242 47796 56252
rect 48972 56308 49028 56318
rect 48972 56214 49028 56252
rect 49980 56308 50036 59200
rect 52220 57428 52276 59200
rect 52220 57372 52388 57428
rect 50556 56476 50820 56486
rect 50612 56420 50660 56476
rect 50716 56420 50764 56476
rect 50556 56410 50820 56420
rect 49980 56242 50036 56252
rect 52220 56308 52276 56318
rect 52220 56214 52276 56252
rect 47740 56084 47796 56094
rect 47964 56084 48020 56094
rect 47740 56082 48020 56084
rect 47740 56030 47742 56082
rect 47794 56030 47966 56082
rect 48018 56030 48020 56082
rect 47740 56028 48020 56030
rect 45500 55346 45556 55356
rect 46732 55412 46788 55422
rect 46732 55318 46788 55356
rect 45724 55298 45780 55310
rect 45724 55246 45726 55298
rect 45778 55246 45780 55298
rect 43484 55074 43764 55076
rect 43484 55022 43598 55074
rect 43650 55022 43764 55074
rect 43484 55020 43764 55022
rect 45388 55076 45444 55086
rect 45724 55076 45780 55246
rect 45388 55074 45780 55076
rect 45388 55022 45390 55074
rect 45442 55022 45780 55074
rect 45388 55020 45780 55022
rect 43484 53956 43540 55020
rect 43596 54982 43652 55020
rect 43484 53890 43540 53900
rect 42476 53620 42532 53630
rect 42476 53618 42644 53620
rect 42476 53566 42478 53618
rect 42530 53566 42644 53618
rect 42476 53564 42644 53566
rect 42476 53554 42532 53564
rect 42252 53508 42308 53518
rect 42252 53506 42420 53508
rect 42252 53454 42254 53506
rect 42306 53454 42420 53506
rect 42252 53452 42420 53454
rect 42252 53442 42308 53452
rect 41692 52334 41694 52386
rect 41746 52334 41748 52386
rect 41244 51492 41300 51502
rect 41020 51438 41022 51490
rect 41074 51438 41076 51490
rect 41020 51380 41076 51438
rect 41020 51314 41076 51324
rect 41132 51436 41244 51492
rect 40908 50708 40964 50718
rect 40908 50614 40964 50652
rect 41020 50036 41076 50046
rect 41132 50036 41188 51436
rect 41244 51398 41300 51436
rect 41244 50708 41300 50718
rect 41468 50708 41524 51772
rect 41692 51716 41748 52334
rect 41916 52668 42084 52724
rect 41916 52162 41972 52668
rect 41916 52110 41918 52162
rect 41970 52110 41972 52162
rect 41916 52098 41972 52110
rect 42252 52052 42308 52062
rect 42252 51958 42308 51996
rect 41580 51660 41748 51716
rect 41580 51156 41636 51660
rect 41804 51604 41860 51614
rect 41580 51062 41636 51100
rect 41692 51602 41860 51604
rect 41692 51550 41806 51602
rect 41858 51550 41860 51602
rect 41692 51548 41860 51550
rect 41692 51044 41748 51548
rect 41804 51538 41860 51548
rect 42252 51604 42308 51614
rect 42364 51604 42420 53452
rect 42588 52836 42644 53564
rect 42700 52948 42756 52958
rect 42700 52854 42756 52892
rect 42588 52612 42644 52780
rect 42588 52556 42756 52612
rect 42700 52274 42756 52556
rect 42700 52222 42702 52274
rect 42754 52222 42756 52274
rect 42700 52210 42756 52222
rect 42588 52164 42644 52174
rect 42308 51548 42420 51604
rect 42476 52162 42644 52164
rect 42476 52110 42590 52162
rect 42642 52110 42644 52162
rect 42476 52108 42644 52110
rect 42252 51510 42308 51548
rect 41804 51378 41860 51390
rect 41804 51326 41806 51378
rect 41858 51326 41860 51378
rect 41804 51268 41860 51326
rect 42140 51268 42196 51278
rect 41804 51266 42196 51268
rect 41804 51214 42142 51266
rect 42194 51214 42196 51266
rect 41804 51212 42196 51214
rect 42140 51202 42196 51212
rect 42476 51154 42532 52108
rect 42588 52098 42644 52108
rect 43036 52164 43092 52174
rect 43148 52164 43204 53676
rect 43036 52162 43204 52164
rect 43036 52110 43038 52162
rect 43090 52110 43204 52162
rect 43036 52108 43204 52110
rect 44604 53844 44660 53854
rect 43036 52098 43092 52108
rect 42476 51102 42478 51154
rect 42530 51102 42532 51154
rect 41692 50988 42084 51044
rect 41300 50652 41524 50708
rect 42028 50706 42084 50988
rect 42028 50654 42030 50706
rect 42082 50654 42084 50706
rect 41244 50594 41300 50652
rect 42028 50642 42084 50654
rect 42476 50708 42532 51102
rect 42476 50642 42532 50652
rect 44156 50708 44212 50718
rect 44156 50614 44212 50652
rect 41244 50542 41246 50594
rect 41298 50542 41300 50594
rect 41244 50530 41300 50542
rect 41020 50034 41188 50036
rect 41020 49982 41022 50034
rect 41074 49982 41188 50034
rect 41020 49980 41188 49982
rect 41020 49970 41076 49980
rect 42700 47460 42756 47470
rect 42700 47366 42756 47404
rect 41244 47348 41300 47358
rect 41132 47012 41188 47022
rect 40908 46900 40964 46910
rect 40908 46786 40964 46844
rect 40908 46734 40910 46786
rect 40962 46734 40964 46786
rect 40908 46722 40964 46734
rect 41132 46786 41188 46956
rect 41244 46898 41300 47292
rect 42028 47348 42084 47358
rect 42028 47254 42084 47292
rect 41244 46846 41246 46898
rect 41298 46846 41300 46898
rect 41244 46834 41300 46846
rect 41132 46734 41134 46786
rect 41186 46734 41188 46786
rect 41132 46722 41188 46734
rect 41468 46788 41524 46798
rect 41524 46732 41972 46788
rect 41468 46694 41524 46732
rect 41020 46004 41076 46014
rect 40796 46002 41636 46004
rect 40796 45950 41022 46002
rect 41074 45950 41636 46002
rect 40796 45948 41636 45950
rect 40236 45780 40292 45790
rect 40236 45330 40292 45724
rect 40236 45278 40238 45330
rect 40290 45278 40292 45330
rect 40236 45266 40292 45278
rect 39676 45054 39678 45106
rect 39730 45054 39732 45106
rect 39676 43652 39732 45054
rect 40124 45106 40180 45118
rect 40124 45054 40126 45106
rect 40178 45054 40180 45106
rect 40124 44996 40180 45054
rect 40124 44930 40180 44940
rect 40348 45108 40404 45118
rect 40348 43708 40404 45052
rect 40796 44548 40852 45948
rect 41020 45938 41076 45948
rect 41580 45890 41636 45948
rect 41580 45838 41582 45890
rect 41634 45838 41636 45890
rect 41580 45826 41636 45838
rect 41916 45890 41972 46732
rect 41916 45838 41918 45890
rect 41970 45838 41972 45890
rect 41916 45826 41972 45838
rect 41356 45780 41412 45790
rect 41356 45686 41412 45724
rect 41804 45666 41860 45678
rect 41804 45614 41806 45666
rect 41858 45614 41860 45666
rect 41804 45332 41860 45614
rect 41804 45276 42420 45332
rect 42364 45218 42420 45276
rect 42364 45166 42366 45218
rect 42418 45166 42420 45218
rect 42364 45154 42420 45166
rect 40796 44482 40852 44492
rect 41580 45106 41636 45118
rect 41580 45054 41582 45106
rect 41634 45054 41636 45106
rect 39676 43586 39732 43596
rect 40236 43652 40404 43708
rect 40796 43652 41300 43708
rect 40012 43540 40068 43550
rect 40012 43446 40068 43484
rect 40236 43428 40292 43652
rect 39564 43148 40180 43204
rect 40124 42754 40180 43148
rect 40124 42702 40126 42754
rect 40178 42702 40180 42754
rect 40124 42690 40180 42702
rect 39452 42590 39454 42642
rect 39506 42590 39508 42642
rect 39452 42578 39508 42590
rect 40236 42644 40292 43372
rect 40796 42754 40852 43652
rect 41244 43650 41300 43652
rect 41244 43598 41246 43650
rect 41298 43598 41300 43650
rect 41244 43586 41300 43598
rect 40796 42702 40798 42754
rect 40850 42702 40852 42754
rect 40796 42690 40852 42702
rect 41020 43540 41076 43550
rect 41020 42756 41076 43484
rect 41132 43538 41188 43550
rect 41132 43486 41134 43538
rect 41186 43486 41188 43538
rect 41132 43428 41188 43486
rect 41132 43362 41188 43372
rect 41356 43538 41412 43550
rect 41356 43486 41358 43538
rect 41410 43486 41412 43538
rect 41356 42868 41412 43486
rect 41580 43540 41636 45054
rect 44492 44996 44548 45006
rect 44492 44902 44548 44940
rect 41580 43474 41636 43484
rect 41692 43652 41748 43662
rect 41692 43538 41748 43596
rect 41692 43486 41694 43538
rect 41746 43486 41748 43538
rect 41692 43474 41748 43486
rect 41244 42812 41356 42868
rect 41132 42756 41188 42766
rect 41020 42754 41188 42756
rect 41020 42702 41134 42754
rect 41186 42702 41188 42754
rect 41020 42700 41188 42702
rect 41132 42690 41188 42700
rect 40236 42578 40292 42588
rect 40460 42644 40516 42654
rect 40460 42530 40516 42588
rect 40460 42478 40462 42530
rect 40514 42478 40516 42530
rect 40460 42466 40516 42478
rect 40572 42642 40628 42654
rect 40572 42590 40574 42642
rect 40626 42590 40628 42642
rect 36988 40402 37044 42364
rect 37772 41972 37828 41982
rect 37772 40514 37828 41916
rect 39900 41860 39956 41870
rect 39900 41766 39956 41804
rect 40460 41860 40516 41870
rect 40572 41860 40628 42590
rect 41020 42084 41076 42094
rect 41244 42084 41300 42812
rect 41356 42802 41412 42812
rect 44044 42868 44100 42878
rect 44044 42774 44100 42812
rect 41916 42644 41972 42654
rect 41916 42550 41972 42588
rect 44604 42420 44660 53788
rect 44828 52836 44884 52846
rect 44828 52742 44884 52780
rect 45388 48916 45444 55020
rect 45388 48850 45444 48860
rect 47740 47572 47796 56028
rect 47964 56018 48020 56028
rect 51212 56082 51268 56094
rect 51212 56030 51214 56082
rect 51266 56030 51268 56082
rect 51212 55468 51268 56030
rect 50876 55412 51268 55468
rect 52332 55412 52388 57372
rect 54460 56308 54516 59200
rect 54460 56242 54516 56252
rect 56028 56308 56084 56318
rect 56028 56214 56084 56252
rect 54572 56084 54628 56094
rect 55020 56084 55076 56094
rect 54572 56082 55076 56084
rect 54572 56030 54574 56082
rect 54626 56030 55022 56082
rect 55074 56030 55076 56082
rect 54572 56028 55076 56030
rect 50876 55074 50932 55412
rect 52332 55346 52388 55356
rect 53676 55412 53732 55422
rect 53676 55318 53732 55356
rect 52668 55298 52724 55310
rect 52668 55246 52670 55298
rect 52722 55246 52724 55298
rect 50876 55022 50878 55074
rect 50930 55022 50932 55074
rect 50556 54908 50820 54918
rect 50612 54852 50660 54908
rect 50716 54852 50764 54908
rect 50556 54842 50820 54852
rect 50876 53844 50932 55022
rect 47740 47506 47796 47516
rect 50316 53788 50932 53844
rect 52108 55076 52164 55086
rect 52668 55076 52724 55246
rect 52108 55074 52724 55076
rect 52108 55022 52110 55074
rect 52162 55022 52724 55074
rect 52108 55020 52724 55022
rect 50316 46004 50372 53788
rect 50556 53340 50820 53350
rect 50612 53284 50660 53340
rect 50716 53284 50764 53340
rect 50556 53274 50820 53284
rect 50556 51772 50820 51782
rect 50612 51716 50660 51772
rect 50716 51716 50764 51772
rect 50556 51706 50820 51716
rect 50556 50204 50820 50214
rect 50612 50148 50660 50204
rect 50716 50148 50764 50204
rect 50556 50138 50820 50148
rect 50556 48636 50820 48646
rect 50612 48580 50660 48636
rect 50716 48580 50764 48636
rect 50556 48570 50820 48580
rect 50556 47068 50820 47078
rect 50612 47012 50660 47068
rect 50716 47012 50764 47068
rect 50556 47002 50820 47012
rect 50316 45938 50372 45948
rect 50556 45500 50820 45510
rect 50612 45444 50660 45500
rect 50716 45444 50764 45500
rect 50556 45434 50820 45444
rect 50556 43932 50820 43942
rect 50612 43876 50660 43932
rect 50716 43876 50764 43932
rect 50556 43866 50820 43876
rect 44604 42354 44660 42364
rect 50556 42364 50820 42374
rect 50612 42308 50660 42364
rect 50716 42308 50764 42364
rect 50556 42298 50820 42308
rect 41020 42082 41300 42084
rect 41020 42030 41022 42082
rect 41074 42030 41300 42082
rect 41020 42028 41300 42030
rect 41020 42018 41076 42028
rect 40516 41804 40628 41860
rect 40460 41794 40516 41804
rect 40908 41746 40964 41758
rect 40908 41694 40910 41746
rect 40962 41694 40964 41746
rect 40908 41188 40964 41694
rect 40908 41122 40964 41132
rect 52108 40964 52164 55020
rect 54572 53844 54628 56028
rect 55020 56018 55076 56028
rect 56700 55410 56756 59200
rect 56700 55358 56702 55410
rect 56754 55358 56756 55410
rect 56700 55346 56756 55358
rect 55580 55298 55636 55310
rect 55580 55246 55582 55298
rect 55634 55246 55636 55298
rect 55244 54404 55300 54414
rect 55580 54404 55636 55246
rect 55244 54402 55636 54404
rect 55244 54350 55246 54402
rect 55298 54350 55636 54402
rect 55244 54348 55636 54350
rect 55244 54338 55300 54348
rect 54572 53778 54628 53788
rect 55356 44436 55412 54348
rect 55356 44370 55412 44380
rect 52108 40898 52164 40908
rect 50556 40796 50820 40806
rect 50612 40740 50660 40796
rect 50716 40740 50764 40796
rect 50556 40730 50820 40740
rect 37772 40462 37774 40514
rect 37826 40462 37828 40514
rect 37772 40450 37828 40462
rect 36988 40350 36990 40402
rect 37042 40350 37044 40402
rect 36428 38612 36708 38668
rect 36764 38834 36820 38846
rect 36764 38782 36766 38834
rect 36818 38782 36820 38834
rect 36428 38162 36484 38612
rect 36428 38110 36430 38162
rect 36482 38110 36484 38162
rect 36428 38052 36484 38110
rect 36428 37986 36484 37996
rect 35868 37326 35870 37378
rect 35922 37326 35924 37378
rect 35868 37314 35924 37326
rect 35644 37202 35700 37212
rect 36204 36484 36260 36494
rect 36764 36484 36820 38782
rect 36988 38724 37044 40350
rect 39900 40290 39956 40302
rect 39900 40238 39902 40290
rect 39954 40238 39956 40290
rect 38220 38948 38276 38958
rect 38220 38854 38276 38892
rect 36988 38658 37044 38668
rect 37436 38834 37492 38846
rect 37436 38782 37438 38834
rect 37490 38782 37492 38834
rect 37436 38724 37492 38782
rect 37436 38658 37492 38668
rect 37212 38276 37268 38286
rect 37212 38162 37268 38220
rect 37772 38276 37828 38286
rect 37772 38182 37828 38220
rect 39340 38276 39396 38286
rect 39900 38276 39956 40238
rect 50556 39228 50820 39238
rect 50612 39172 50660 39228
rect 50716 39172 50764 39228
rect 50556 39162 50820 39172
rect 40348 38724 40404 38734
rect 39396 38220 39508 38276
rect 39340 38210 39396 38220
rect 37212 38110 37214 38162
rect 37266 38110 37268 38162
rect 37212 38098 37268 38110
rect 37996 38050 38052 38062
rect 38220 38052 38276 38062
rect 37996 37998 37998 38050
rect 38050 37998 38052 38050
rect 37996 37156 38052 37998
rect 37996 37062 38052 37100
rect 38108 38050 38276 38052
rect 38108 37998 38222 38050
rect 38274 37998 38276 38050
rect 38108 37996 38276 37998
rect 38108 37380 38164 37996
rect 38220 37986 38276 37996
rect 38444 38052 38500 38062
rect 36204 36482 36820 36484
rect 36204 36430 36206 36482
rect 36258 36430 36820 36482
rect 36204 36428 36820 36430
rect 37324 36594 37380 36606
rect 37324 36542 37326 36594
rect 37378 36542 37380 36594
rect 35532 35858 35588 35868
rect 35644 36370 35700 36382
rect 35644 36318 35646 36370
rect 35698 36318 35700 36370
rect 35644 35812 35700 36318
rect 34748 35410 34804 35420
rect 34972 35700 35028 35710
rect 34524 34748 34692 34804
rect 34860 34802 34916 34814
rect 34860 34750 34862 34802
rect 34914 34750 34916 34802
rect 34524 32676 34580 34748
rect 34748 32900 34804 32910
rect 34524 32610 34580 32620
rect 34636 32844 34748 32900
rect 34636 32562 34692 32844
rect 34748 32834 34804 32844
rect 34636 32510 34638 32562
rect 34690 32510 34692 32562
rect 34636 32498 34692 32510
rect 34748 32564 34804 32574
rect 34412 31042 34468 31052
rect 34748 30994 34804 32508
rect 34748 30942 34750 30994
rect 34802 30942 34804 30994
rect 34748 30930 34804 30942
rect 34300 30828 34580 30884
rect 34524 30322 34580 30828
rect 34524 30270 34526 30322
rect 34578 30270 34580 30322
rect 34524 30258 34580 30270
rect 34860 30212 34916 34750
rect 34972 32900 35028 35644
rect 35196 35308 35460 35318
rect 35252 35252 35300 35308
rect 35356 35252 35404 35308
rect 35196 35242 35460 35252
rect 35532 35140 35588 35150
rect 35644 35140 35700 35756
rect 36204 35700 36260 36428
rect 36428 35924 36484 35934
rect 36428 35810 36484 35868
rect 36428 35758 36430 35810
rect 36482 35758 36484 35810
rect 36428 35746 36484 35758
rect 36204 35634 36260 35644
rect 37100 35700 37156 35710
rect 37100 35606 37156 35644
rect 35588 35084 35700 35140
rect 35532 35074 35588 35084
rect 35420 34914 35476 34926
rect 35420 34862 35422 34914
rect 35474 34862 35476 34914
rect 35308 34692 35364 34702
rect 35308 34598 35364 34636
rect 35420 34132 35476 34862
rect 35644 34242 35700 35084
rect 36316 35476 36372 35486
rect 36316 34804 36372 35420
rect 36316 34710 36372 34748
rect 36428 35364 36484 35374
rect 36428 34914 36484 35308
rect 36428 34862 36430 34914
rect 36482 34862 36484 34914
rect 36428 34580 36484 34862
rect 35644 34190 35646 34242
rect 35698 34190 35700 34242
rect 35644 34178 35700 34190
rect 36204 34524 36484 34580
rect 36876 34916 36932 34926
rect 35420 34066 35476 34076
rect 36092 34132 36148 34142
rect 35196 33740 35460 33750
rect 35252 33684 35300 33740
rect 35356 33684 35404 33740
rect 35196 33674 35460 33684
rect 36092 33684 36148 34076
rect 36092 33618 36148 33628
rect 34972 32834 35028 32844
rect 35196 33346 35252 33358
rect 35196 33294 35198 33346
rect 35250 33294 35252 33346
rect 35196 32564 35252 33294
rect 36204 33346 36260 34524
rect 36428 34132 36484 34142
rect 36428 34038 36484 34076
rect 36204 33294 36206 33346
rect 36258 33294 36260 33346
rect 36204 33282 36260 33294
rect 36540 34018 36596 34030
rect 36540 33966 36542 34018
rect 36594 33966 36596 34018
rect 35196 32470 35252 32508
rect 35644 33236 35700 33246
rect 35644 32674 35700 33180
rect 36428 33122 36484 33134
rect 36428 33070 36430 33122
rect 36482 33070 36484 33122
rect 36428 32900 36484 33070
rect 36428 32834 36484 32844
rect 35644 32622 35646 32674
rect 35698 32622 35700 32674
rect 35196 32172 35460 32182
rect 35252 32116 35300 32172
rect 35356 32116 35404 32172
rect 35196 32106 35460 32116
rect 35196 31668 35252 31678
rect 35196 31574 35252 31612
rect 35644 31668 35700 32622
rect 35644 31602 35700 31612
rect 35756 31108 35812 31118
rect 35756 31014 35812 31052
rect 35980 30996 36036 31006
rect 35868 30940 35980 30996
rect 35196 30604 35460 30614
rect 35252 30548 35300 30604
rect 35356 30548 35404 30604
rect 35196 30538 35460 30548
rect 34972 30212 35028 30222
rect 34860 30156 34972 30212
rect 34972 30118 35028 30156
rect 35644 30212 35700 30222
rect 35644 30118 35700 30156
rect 35756 29650 35812 29662
rect 35756 29598 35758 29650
rect 35810 29598 35812 29650
rect 34300 29540 34356 29550
rect 34188 29538 34356 29540
rect 34188 29486 34302 29538
rect 34354 29486 34356 29538
rect 34188 29484 34356 29486
rect 34300 29474 34356 29484
rect 35196 29036 35460 29046
rect 35252 28980 35300 29036
rect 35356 28980 35404 29036
rect 35196 28970 35460 28980
rect 35756 28084 35812 29598
rect 35868 29426 35924 30940
rect 35980 30930 36036 30940
rect 36540 30436 36596 33966
rect 36876 30996 36932 34860
rect 37100 34804 37156 34814
rect 37100 34710 37156 34748
rect 37212 34692 37268 34702
rect 37212 34598 37268 34636
rect 37324 33684 37380 36542
rect 37996 36484 38052 36494
rect 38108 36484 38164 37324
rect 38052 36428 38164 36484
rect 37996 36390 38052 36428
rect 38444 36036 38500 37996
rect 38668 37266 38724 37278
rect 38668 37214 38670 37266
rect 38722 37214 38724 37266
rect 38668 37156 38724 37214
rect 38108 35980 38444 36036
rect 37436 35812 37492 35822
rect 37436 35718 37492 35756
rect 37660 35810 37716 35822
rect 37660 35758 37662 35810
rect 37714 35758 37716 35810
rect 37660 34804 37716 35758
rect 37660 34738 37716 34748
rect 37324 33618 37380 33628
rect 37100 33348 37156 33358
rect 37100 33254 37156 33292
rect 37212 33124 37268 33134
rect 37212 33030 37268 33068
rect 37660 33122 37716 33134
rect 37660 33070 37662 33122
rect 37714 33070 37716 33122
rect 37660 32788 37716 33070
rect 37660 32722 37716 32732
rect 37324 32676 37380 32686
rect 37324 32582 37380 32620
rect 36876 30902 36932 30940
rect 36988 31666 37044 31678
rect 36988 31614 36990 31666
rect 37042 31614 37044 31666
rect 36428 30380 36596 30436
rect 35980 30100 36036 30110
rect 35980 30006 36036 30044
rect 35868 29374 35870 29426
rect 35922 29374 35924 29426
rect 35868 29362 35924 29374
rect 35756 28018 35812 28028
rect 35196 27468 35460 27478
rect 35252 27412 35300 27468
rect 35356 27412 35404 27468
rect 35196 27402 35460 27412
rect 30492 26852 30772 26908
rect 32060 26852 32228 26908
rect 33628 26852 34132 26908
rect 28252 26628 28308 26638
rect 28252 25618 28308 26572
rect 28252 25566 28254 25618
rect 28306 25566 28308 25618
rect 28252 25554 28308 25566
rect 29260 25284 29316 25294
rect 29260 25190 29316 25228
rect 30492 24836 30548 26852
rect 32060 24948 32116 26852
rect 33628 25620 33684 26852
rect 35196 25900 35460 25910
rect 35252 25844 35300 25900
rect 35356 25844 35404 25900
rect 35196 25834 35460 25844
rect 33628 25554 33684 25564
rect 36428 25284 36484 30380
rect 36988 30212 37044 31614
rect 37436 31668 37492 31678
rect 37212 31556 37268 31566
rect 37212 31462 37268 31500
rect 37436 30882 37492 31612
rect 37436 30830 37438 30882
rect 37490 30830 37492 30882
rect 36988 30146 37044 30156
rect 37212 30212 37268 30222
rect 37212 30118 37268 30156
rect 36540 30100 36596 30110
rect 36540 30006 36596 30044
rect 37436 29538 37492 30830
rect 38108 30996 38164 35980
rect 38444 35970 38500 35980
rect 38556 36484 38612 36494
rect 38668 36484 38724 37100
rect 38556 36482 38724 36484
rect 38556 36430 38558 36482
rect 38610 36430 38724 36482
rect 38556 36428 38724 36430
rect 39116 37154 39172 37166
rect 39116 37102 39118 37154
rect 39170 37102 39172 37154
rect 38556 35698 38612 36428
rect 38556 35646 38558 35698
rect 38610 35646 38612 35698
rect 38556 35634 38612 35646
rect 39004 36260 39060 36270
rect 39004 35700 39060 36204
rect 38668 35140 38724 35150
rect 38556 35084 38668 35140
rect 38556 34916 38612 35084
rect 38668 35074 38724 35084
rect 38556 34822 38612 34860
rect 39004 34914 39060 35644
rect 39004 34862 39006 34914
rect 39058 34862 39060 34914
rect 39004 34850 39060 34862
rect 39116 35364 39172 37102
rect 39340 36594 39396 36606
rect 39340 36542 39342 36594
rect 39394 36542 39396 36594
rect 39228 35924 39284 35934
rect 39228 35810 39284 35868
rect 39228 35758 39230 35810
rect 39282 35758 39284 35810
rect 39228 35746 39284 35758
rect 38892 34018 38948 34030
rect 38892 33966 38894 34018
rect 38946 33966 38948 34018
rect 38220 33684 38276 33694
rect 38220 31780 38276 33628
rect 38892 33684 38948 33966
rect 38892 33618 38948 33628
rect 39116 33460 39172 35308
rect 39340 35140 39396 36542
rect 39340 35074 39396 35084
rect 38444 33404 39172 33460
rect 38444 32562 38500 33404
rect 39116 33346 39172 33404
rect 39116 33294 39118 33346
rect 39170 33294 39172 33346
rect 39116 33282 39172 33294
rect 39452 34130 39508 38220
rect 39900 38210 39956 38220
rect 40236 38722 40404 38724
rect 40236 38670 40350 38722
rect 40402 38670 40404 38722
rect 40236 38668 40404 38670
rect 39900 37492 39956 37502
rect 40236 37492 40292 38668
rect 40348 38658 40404 38668
rect 50556 37660 50820 37670
rect 50612 37604 50660 37660
rect 50716 37604 50764 37660
rect 50556 37594 50820 37604
rect 39900 37490 40292 37492
rect 39900 37438 39902 37490
rect 39954 37438 40292 37490
rect 39900 37436 40292 37438
rect 39900 37426 39956 37436
rect 39564 37380 39620 37390
rect 39564 37286 39620 37324
rect 40236 37378 40292 37436
rect 40236 37326 40238 37378
rect 40290 37326 40292 37378
rect 40236 37314 40292 37326
rect 40348 37042 40404 37054
rect 40348 36990 40350 37042
rect 40402 36990 40404 37042
rect 40124 36260 40180 36270
rect 40348 36260 40404 36990
rect 40908 36260 40964 36270
rect 40348 36258 41076 36260
rect 40348 36206 40910 36258
rect 40962 36206 41076 36258
rect 40348 36204 41076 36206
rect 40124 36166 40180 36204
rect 40908 36194 40964 36204
rect 40348 36036 40404 36046
rect 40348 35922 40404 35980
rect 40348 35870 40350 35922
rect 40402 35870 40404 35922
rect 40348 35858 40404 35870
rect 40908 36036 40964 36046
rect 40908 35922 40964 35980
rect 40908 35870 40910 35922
rect 40962 35870 40964 35922
rect 40908 35858 40964 35870
rect 39676 35698 39732 35710
rect 39676 35646 39678 35698
rect 39730 35646 39732 35698
rect 39676 35588 39732 35646
rect 39452 34078 39454 34130
rect 39506 34078 39508 34130
rect 39452 33348 39508 34078
rect 39564 34804 39620 34814
rect 39676 34804 39732 35532
rect 39564 34802 39732 34804
rect 39564 34750 39566 34802
rect 39618 34750 39732 34802
rect 39564 34748 39732 34750
rect 39564 34132 39620 34748
rect 39564 34066 39620 34076
rect 40124 34132 40180 34142
rect 39452 33282 39508 33292
rect 39676 33572 39732 33582
rect 38444 32510 38446 32562
rect 38498 32510 38500 32562
rect 38444 32498 38500 32510
rect 38668 33234 38724 33246
rect 38668 33182 38670 33234
rect 38722 33182 38724 33234
rect 38668 33124 38724 33182
rect 38668 32564 38724 33068
rect 39116 32900 39172 32910
rect 38780 32564 38836 32574
rect 38668 32562 38836 32564
rect 38668 32510 38782 32562
rect 38834 32510 38836 32562
rect 38668 32508 38836 32510
rect 38780 32498 38836 32508
rect 38668 31780 38724 31790
rect 38220 31778 38724 31780
rect 38220 31726 38670 31778
rect 38722 31726 38724 31778
rect 38220 31724 38724 31726
rect 38220 30996 38276 31006
rect 38108 30994 38276 30996
rect 38108 30942 38222 30994
rect 38274 30942 38276 30994
rect 38108 30940 38276 30942
rect 38108 30212 38164 30940
rect 38220 30930 38276 30940
rect 38108 30146 38164 30156
rect 37436 29486 37438 29538
rect 37490 29486 37492 29538
rect 37436 29474 37492 29486
rect 38108 29428 38164 29438
rect 38444 29428 38500 31724
rect 38668 31714 38724 31724
rect 39116 31778 39172 32844
rect 39116 31726 39118 31778
rect 39170 31726 39172 31778
rect 39116 31714 39172 31726
rect 39452 32450 39508 32462
rect 39452 32398 39454 32450
rect 39506 32398 39508 32450
rect 39452 31108 39508 32398
rect 39676 31666 39732 33516
rect 40124 33234 40180 34076
rect 40124 33182 40126 33234
rect 40178 33182 40180 33234
rect 40124 33170 40180 33182
rect 40908 33348 40964 33358
rect 41020 33348 41076 36204
rect 50556 36092 50820 36102
rect 50612 36036 50660 36092
rect 50716 36036 50764 36092
rect 50556 36026 50820 36036
rect 41356 35588 41412 35598
rect 41356 35494 41412 35532
rect 41468 34804 41524 34814
rect 41244 33348 41300 33358
rect 41020 33346 41300 33348
rect 41020 33294 41246 33346
rect 41298 33294 41300 33346
rect 41020 33292 41300 33294
rect 40908 32786 40964 33292
rect 41244 33282 41300 33292
rect 40908 32734 40910 32786
rect 40962 32734 40964 32786
rect 40908 32722 40964 32734
rect 41468 32674 41524 34748
rect 50556 34524 50820 34534
rect 50612 34468 50660 34524
rect 50716 34468 50764 34524
rect 50556 34458 50820 34468
rect 50556 32956 50820 32966
rect 50612 32900 50660 32956
rect 50716 32900 50764 32956
rect 50556 32890 50820 32900
rect 41468 32622 41470 32674
rect 41522 32622 41524 32674
rect 41468 32610 41524 32622
rect 39676 31614 39678 31666
rect 39730 31614 39732 31666
rect 39676 31602 39732 31614
rect 50556 31388 50820 31398
rect 50612 31332 50660 31388
rect 50716 31332 50764 31388
rect 50556 31322 50820 31332
rect 39452 31042 39508 31052
rect 50556 29820 50820 29830
rect 50612 29764 50660 29820
rect 50716 29764 50764 29820
rect 50556 29754 50820 29764
rect 38108 29426 38500 29428
rect 38108 29374 38110 29426
rect 38162 29374 38500 29426
rect 38108 29372 38500 29374
rect 38108 29362 38164 29372
rect 50556 28252 50820 28262
rect 50612 28196 50660 28252
rect 50716 28196 50764 28252
rect 50556 28186 50820 28196
rect 50556 26684 50820 26694
rect 50612 26628 50660 26684
rect 50716 26628 50764 26684
rect 50556 26618 50820 26628
rect 36428 25218 36484 25228
rect 50556 25116 50820 25126
rect 50612 25060 50660 25116
rect 50716 25060 50764 25116
rect 50556 25050 50820 25060
rect 32060 24882 32116 24892
rect 30492 24770 30548 24780
rect 35196 24332 35460 24342
rect 35252 24276 35300 24332
rect 35356 24276 35404 24332
rect 35196 24266 35460 24276
rect 50556 23548 50820 23558
rect 50612 23492 50660 23548
rect 50716 23492 50764 23548
rect 50556 23482 50820 23492
rect 27916 22866 27972 22876
rect 35196 22764 35460 22774
rect 35252 22708 35300 22764
rect 35356 22708 35404 22764
rect 35196 22698 35460 22708
rect 27804 22642 27860 22652
rect 15596 22482 15988 22484
rect 15596 22430 15598 22482
rect 15650 22430 15988 22482
rect 15596 22428 15988 22430
rect 15596 22418 15652 22428
rect 19836 21980 20100 21990
rect 19892 21924 19940 21980
rect 19996 21924 20044 21980
rect 19836 21914 20100 21924
rect 50556 21980 50820 21990
rect 50612 21924 50660 21980
rect 50716 21924 50764 21980
rect 50556 21914 50820 21924
rect 12684 21634 12740 21644
rect 35196 21196 35460 21206
rect 35252 21140 35300 21196
rect 35356 21140 35404 21196
rect 35196 21130 35460 21140
rect 19836 20412 20100 20422
rect 19892 20356 19940 20412
rect 19996 20356 20044 20412
rect 19836 20346 20100 20356
rect 50556 20412 50820 20422
rect 50612 20356 50660 20412
rect 50716 20356 50764 20412
rect 50556 20346 50820 20356
rect 8092 20132 8260 20188
rect 6524 9986 6580 9996
rect 2492 9602 2548 9614
rect 2492 9550 2494 9602
rect 2546 9550 2548 9602
rect 2492 9268 2548 9550
rect 2492 9202 2548 9212
rect 4476 8652 4740 8662
rect 4532 8596 4580 8652
rect 4636 8596 4684 8652
rect 4476 8586 4740 8596
rect 2492 8036 2548 8046
rect 2492 7942 2548 7980
rect 4476 7084 4740 7094
rect 4532 7028 4580 7084
rect 4636 7028 4684 7084
rect 4476 7018 4740 7028
rect 4476 5516 4740 5526
rect 4532 5460 4580 5516
rect 4636 5460 4684 5516
rect 4476 5450 4740 5460
rect 8204 4564 8260 20132
rect 35196 19628 35460 19638
rect 35252 19572 35300 19628
rect 35356 19572 35404 19628
rect 35196 19562 35460 19572
rect 19836 18844 20100 18854
rect 19892 18788 19940 18844
rect 19996 18788 20044 18844
rect 19836 18778 20100 18788
rect 50556 18844 50820 18854
rect 50612 18788 50660 18844
rect 50716 18788 50764 18844
rect 50556 18778 50820 18788
rect 35196 18060 35460 18070
rect 35252 18004 35300 18060
rect 35356 18004 35404 18060
rect 35196 17994 35460 18004
rect 19836 17276 20100 17286
rect 19892 17220 19940 17276
rect 19996 17220 20044 17276
rect 19836 17210 20100 17220
rect 50556 17276 50820 17286
rect 50612 17220 50660 17276
rect 50716 17220 50764 17276
rect 50556 17210 50820 17220
rect 35196 16492 35460 16502
rect 35252 16436 35300 16492
rect 35356 16436 35404 16492
rect 35196 16426 35460 16436
rect 19836 15708 20100 15718
rect 19892 15652 19940 15708
rect 19996 15652 20044 15708
rect 19836 15642 20100 15652
rect 50556 15708 50820 15718
rect 50612 15652 50660 15708
rect 50716 15652 50764 15708
rect 50556 15642 50820 15652
rect 35196 14924 35460 14934
rect 35252 14868 35300 14924
rect 35356 14868 35404 14924
rect 35196 14858 35460 14868
rect 19836 14140 20100 14150
rect 19892 14084 19940 14140
rect 19996 14084 20044 14140
rect 19836 14074 20100 14084
rect 50556 14140 50820 14150
rect 50612 14084 50660 14140
rect 50716 14084 50764 14140
rect 50556 14074 50820 14084
rect 35196 13356 35460 13366
rect 35252 13300 35300 13356
rect 35356 13300 35404 13356
rect 35196 13290 35460 13300
rect 19836 12572 20100 12582
rect 19892 12516 19940 12572
rect 19996 12516 20044 12572
rect 19836 12506 20100 12516
rect 50556 12572 50820 12582
rect 50612 12516 50660 12572
rect 50716 12516 50764 12572
rect 50556 12506 50820 12516
rect 35196 11788 35460 11798
rect 35252 11732 35300 11788
rect 35356 11732 35404 11788
rect 35196 11722 35460 11732
rect 19836 11004 20100 11014
rect 19892 10948 19940 11004
rect 19996 10948 20044 11004
rect 19836 10938 20100 10948
rect 50556 11004 50820 11014
rect 50612 10948 50660 11004
rect 50716 10948 50764 11004
rect 50556 10938 50820 10948
rect 35196 10220 35460 10230
rect 35252 10164 35300 10220
rect 35356 10164 35404 10220
rect 35196 10154 35460 10164
rect 19836 9436 20100 9446
rect 19892 9380 19940 9436
rect 19996 9380 20044 9436
rect 19836 9370 20100 9380
rect 50556 9436 50820 9446
rect 50612 9380 50660 9436
rect 50716 9380 50764 9436
rect 50556 9370 50820 9380
rect 35196 8652 35460 8662
rect 35252 8596 35300 8652
rect 35356 8596 35404 8652
rect 35196 8586 35460 8596
rect 19836 7868 20100 7878
rect 19892 7812 19940 7868
rect 19996 7812 20044 7868
rect 19836 7802 20100 7812
rect 50556 7868 50820 7878
rect 50612 7812 50660 7868
rect 50716 7812 50764 7868
rect 50556 7802 50820 7812
rect 35196 7084 35460 7094
rect 35252 7028 35300 7084
rect 35356 7028 35404 7084
rect 35196 7018 35460 7028
rect 19836 6300 20100 6310
rect 19892 6244 19940 6300
rect 19996 6244 20044 6300
rect 19836 6234 20100 6244
rect 50556 6300 50820 6310
rect 50612 6244 50660 6300
rect 50716 6244 50764 6300
rect 50556 6234 50820 6244
rect 35196 5516 35460 5526
rect 35252 5460 35300 5516
rect 35356 5460 35404 5516
rect 35196 5450 35460 5460
rect 19836 4732 20100 4742
rect 19892 4676 19940 4732
rect 19996 4676 20044 4732
rect 19836 4666 20100 4676
rect 50556 4732 50820 4742
rect 50612 4676 50660 4732
rect 50716 4676 50764 4732
rect 50556 4666 50820 4676
rect 8204 4498 8260 4508
rect 2492 4226 2548 4238
rect 2492 4174 2494 4226
rect 2546 4174 2548 4226
rect 2492 3892 2548 4174
rect 4476 3948 4740 3958
rect 4532 3892 4580 3948
rect 4636 3892 4684 3948
rect 4476 3882 4740 3892
rect 35196 3948 35460 3958
rect 35252 3892 35300 3948
rect 35356 3892 35404 3948
rect 35196 3882 35460 3892
rect 2492 3826 2548 3836
rect 2268 3666 2436 3668
rect 2268 3614 2270 3666
rect 2322 3614 2436 3666
rect 2268 3612 2436 3614
rect 2268 3602 2324 3612
rect 1708 3442 1764 3454
rect 1708 3390 1710 3442
rect 1762 3390 1764 3442
rect 1708 3332 1764 3390
rect 1708 2100 1764 3276
rect 2716 3442 2772 3454
rect 2716 3390 2718 3442
rect 2770 3390 2772 3442
rect 2716 3332 2772 3390
rect 2716 3266 2772 3276
rect 19836 3164 20100 3174
rect 19892 3108 19940 3164
rect 19996 3108 20044 3164
rect 19836 3098 20100 3108
rect 50556 3164 50820 3174
rect 50612 3108 50660 3164
rect 50716 3108 50764 3164
rect 50556 3098 50820 3108
rect 1708 2034 1764 2044
<< via2 >>
rect 2156 57596 2212 57652
rect 1708 55804 1764 55860
rect 2156 56028 2212 56084
rect 1372 54572 1428 54628
rect 1148 39564 1204 39620
rect 1036 35756 1092 35812
rect 1708 54012 1764 54068
rect 1708 52780 1764 52836
rect 1708 52220 1764 52276
rect 1820 51212 1876 51268
rect 1708 50706 1764 50708
rect 1708 50654 1710 50706
rect 1710 50654 1762 50706
rect 1762 50654 1764 50706
rect 1708 50652 1764 50654
rect 1708 50428 1764 50484
rect 2604 56082 2660 56084
rect 2604 56030 2606 56082
rect 2606 56030 2658 56082
rect 2658 56030 2660 56082
rect 2604 56028 2660 56030
rect 2044 54626 2100 54628
rect 2044 54574 2046 54626
rect 2046 54574 2098 54626
rect 2098 54574 2100 54626
rect 2044 54572 2100 54574
rect 2492 54012 2548 54068
rect 2044 51490 2100 51492
rect 2044 51438 2046 51490
rect 2046 51438 2098 51490
rect 2098 51438 2100 51490
rect 2044 51436 2100 51438
rect 2492 52834 2548 52836
rect 2492 52782 2494 52834
rect 2494 52782 2546 52834
rect 2546 52782 2548 52834
rect 2492 52780 2548 52782
rect 2492 51266 2548 51268
rect 2492 51214 2494 51266
rect 2494 51214 2546 51266
rect 2546 51214 2548 51266
rect 2492 51212 2548 51214
rect 1708 48636 1764 48692
rect 1708 46844 1764 46900
rect 1708 45052 1764 45108
rect 1372 36316 1428 36372
rect 1484 44828 1540 44884
rect 1148 29708 1204 29764
rect 1260 32396 1316 32452
rect 1036 23436 1092 23492
rect 1148 26908 1204 26964
rect 1148 15148 1204 15204
rect 2156 47628 2212 47684
rect 2492 48636 2548 48692
rect 3164 55804 3220 55860
rect 4476 55690 4532 55692
rect 4476 55638 4478 55690
rect 4478 55638 4530 55690
rect 4530 55638 4532 55690
rect 4476 55636 4532 55638
rect 4580 55690 4636 55692
rect 4580 55638 4582 55690
rect 4582 55638 4634 55690
rect 4634 55638 4636 55690
rect 4580 55636 4636 55638
rect 4684 55690 4740 55692
rect 4684 55638 4686 55690
rect 4686 55638 4738 55690
rect 4738 55638 4740 55690
rect 4684 55636 4740 55638
rect 19836 56474 19892 56476
rect 19836 56422 19838 56474
rect 19838 56422 19890 56474
rect 19890 56422 19892 56474
rect 19836 56420 19892 56422
rect 19940 56474 19996 56476
rect 19940 56422 19942 56474
rect 19942 56422 19994 56474
rect 19994 56422 19996 56474
rect 19940 56420 19996 56422
rect 20044 56474 20100 56476
rect 20044 56422 20046 56474
rect 20046 56422 20098 56474
rect 20098 56422 20100 56474
rect 20044 56420 20100 56422
rect 5852 55132 5908 55188
rect 4476 54122 4532 54124
rect 4476 54070 4478 54122
rect 4478 54070 4530 54122
rect 4530 54070 4532 54122
rect 4476 54068 4532 54070
rect 4580 54122 4636 54124
rect 4580 54070 4582 54122
rect 4582 54070 4634 54122
rect 4634 54070 4636 54122
rect 4580 54068 4636 54070
rect 4684 54122 4740 54124
rect 4684 54070 4686 54122
rect 4686 54070 4738 54122
rect 4738 54070 4740 54122
rect 4684 54068 4740 54070
rect 2940 53788 2996 53844
rect 5740 53788 5796 53844
rect 4476 52554 4532 52556
rect 4476 52502 4478 52554
rect 4478 52502 4530 52554
rect 4530 52502 4532 52554
rect 4476 52500 4532 52502
rect 4580 52554 4636 52556
rect 4580 52502 4582 52554
rect 4582 52502 4634 52554
rect 4634 52502 4636 52554
rect 4580 52500 4636 52502
rect 4684 52554 4740 52556
rect 4684 52502 4686 52554
rect 4686 52502 4738 52554
rect 4738 52502 4740 52554
rect 4684 52500 4740 52502
rect 3836 51884 3892 51940
rect 2716 51436 2772 51492
rect 3276 50652 3332 50708
rect 2492 47404 2548 47460
rect 1820 43260 1876 43316
rect 2044 43596 2100 43652
rect 2044 43372 2100 43428
rect 2492 46898 2548 46900
rect 2492 46846 2494 46898
rect 2494 46846 2546 46898
rect 2546 46846 2548 46898
rect 2492 46844 2548 46846
rect 2268 45052 2324 45108
rect 2492 45106 2548 45108
rect 2492 45054 2494 45106
rect 2494 45054 2546 45106
rect 2546 45054 2548 45106
rect 2492 45052 2548 45054
rect 2268 44044 2324 44100
rect 4396 51378 4452 51380
rect 4396 51326 4398 51378
rect 4398 51326 4450 51378
rect 4450 51326 4452 51378
rect 4396 51324 4452 51326
rect 5180 51324 5236 51380
rect 5068 51266 5124 51268
rect 5068 51214 5070 51266
rect 5070 51214 5122 51266
rect 5122 51214 5124 51266
rect 5068 51212 5124 51214
rect 4476 50986 4532 50988
rect 4476 50934 4478 50986
rect 4478 50934 4530 50986
rect 4530 50934 4532 50986
rect 4476 50932 4532 50934
rect 4580 50986 4636 50988
rect 4580 50934 4582 50986
rect 4582 50934 4634 50986
rect 4634 50934 4636 50986
rect 4580 50932 4636 50934
rect 4684 50986 4740 50988
rect 4684 50934 4686 50986
rect 4686 50934 4738 50986
rect 4738 50934 4740 50986
rect 4684 50932 4740 50934
rect 3836 49922 3892 49924
rect 3836 49870 3838 49922
rect 3838 49870 3890 49922
rect 3890 49870 3892 49922
rect 3836 49868 3892 49870
rect 4476 49418 4532 49420
rect 4476 49366 4478 49418
rect 4478 49366 4530 49418
rect 4530 49366 4532 49418
rect 4476 49364 4532 49366
rect 4580 49418 4636 49420
rect 4580 49366 4582 49418
rect 4582 49366 4634 49418
rect 4634 49366 4636 49418
rect 4580 49364 4636 49366
rect 4684 49418 4740 49420
rect 4684 49366 4686 49418
rect 4686 49366 4738 49418
rect 4738 49366 4740 49418
rect 4684 49364 4740 49366
rect 3276 47682 3332 47684
rect 3276 47630 3278 47682
rect 3278 47630 3330 47682
rect 3330 47630 3332 47682
rect 3276 47628 3332 47630
rect 3948 47458 4004 47460
rect 3948 47406 3950 47458
rect 3950 47406 4002 47458
rect 4002 47406 4004 47458
rect 3948 47404 4004 47406
rect 2716 44044 2772 44100
rect 2380 43484 2436 43540
rect 1708 41468 1764 41524
rect 1708 40236 1764 40292
rect 1708 39676 1764 39732
rect 1708 37938 1764 37940
rect 1708 37886 1710 37938
rect 1710 37886 1762 37938
rect 1762 37886 1764 37938
rect 1708 37884 1764 37886
rect 2044 41916 2100 41972
rect 2044 39564 2100 39620
rect 3052 45106 3108 45108
rect 3052 45054 3054 45106
rect 3054 45054 3106 45106
rect 3106 45054 3108 45106
rect 3052 45052 3108 45054
rect 3164 44882 3220 44884
rect 3164 44830 3166 44882
rect 3166 44830 3218 44882
rect 3218 44830 3220 44882
rect 3164 44828 3220 44830
rect 2716 43650 2772 43652
rect 2716 43598 2718 43650
rect 2718 43598 2770 43650
rect 2770 43598 2772 43650
rect 2716 43596 2772 43598
rect 2716 42252 2772 42308
rect 2716 41970 2772 41972
rect 2716 41918 2718 41970
rect 2718 41918 2770 41970
rect 2770 41918 2772 41970
rect 2716 41916 2772 41918
rect 3052 42530 3108 42532
rect 3052 42478 3054 42530
rect 3054 42478 3106 42530
rect 3106 42478 3108 42530
rect 3052 42476 3108 42478
rect 3052 42252 3108 42308
rect 2604 41132 2660 41188
rect 2492 41020 2548 41076
rect 2716 41074 2772 41076
rect 2716 41022 2718 41074
rect 2718 41022 2770 41074
rect 2770 41022 2772 41074
rect 2716 41020 2772 41022
rect 3724 47068 3780 47124
rect 4476 47850 4532 47852
rect 4476 47798 4478 47850
rect 4478 47798 4530 47850
rect 4530 47798 4532 47850
rect 4476 47796 4532 47798
rect 4580 47850 4636 47852
rect 4580 47798 4582 47850
rect 4582 47798 4634 47850
rect 4634 47798 4636 47850
rect 4580 47796 4636 47798
rect 4684 47850 4740 47852
rect 4684 47798 4686 47850
rect 4686 47798 4738 47850
rect 4738 47798 4740 47850
rect 4684 47796 4740 47798
rect 4060 47068 4116 47124
rect 7980 52946 8036 52948
rect 7980 52894 7982 52946
rect 7982 52894 8034 52946
rect 8034 52894 8036 52946
rect 7980 52892 8036 52894
rect 7644 51378 7700 51380
rect 7644 51326 7646 51378
rect 7646 51326 7698 51378
rect 7698 51326 7700 51378
rect 7644 51324 7700 51326
rect 5852 50764 5908 50820
rect 7308 50818 7364 50820
rect 7308 50766 7310 50818
rect 7310 50766 7362 50818
rect 7362 50766 7364 50818
rect 7308 50764 7364 50766
rect 5740 47180 5796 47236
rect 6076 48188 6132 48244
rect 4508 46844 4564 46900
rect 4844 46786 4900 46788
rect 4844 46734 4846 46786
rect 4846 46734 4898 46786
rect 4898 46734 4900 46786
rect 4844 46732 4900 46734
rect 4476 46282 4532 46284
rect 4476 46230 4478 46282
rect 4478 46230 4530 46282
rect 4530 46230 4532 46282
rect 4476 46228 4532 46230
rect 4580 46282 4636 46284
rect 4580 46230 4582 46282
rect 4582 46230 4634 46282
rect 4634 46230 4636 46282
rect 4580 46228 4636 46230
rect 4684 46282 4740 46284
rect 4684 46230 4686 46282
rect 4686 46230 4738 46282
rect 4738 46230 4740 46282
rect 4684 46228 4740 46230
rect 4508 45778 4564 45780
rect 4508 45726 4510 45778
rect 4510 45726 4562 45778
rect 4562 45726 4564 45778
rect 4508 45724 4564 45726
rect 4172 45388 4228 45444
rect 4060 45276 4116 45332
rect 3612 43596 3668 43652
rect 3724 43260 3780 43316
rect 2492 40236 2548 40292
rect 2604 39564 2660 39620
rect 1932 37436 1988 37492
rect 1708 37100 1764 37156
rect 1708 36092 1764 36148
rect 2044 36428 2100 36484
rect 1932 36370 1988 36372
rect 1932 36318 1934 36370
rect 1934 36318 1986 36370
rect 1986 36318 1988 36370
rect 1932 36316 1988 36318
rect 1708 34354 1764 34356
rect 1708 34302 1710 34354
rect 1710 34302 1762 34354
rect 1762 34302 1764 34354
rect 1708 34300 1764 34302
rect 1708 33234 1764 33236
rect 1708 33182 1710 33234
rect 1710 33182 1762 33234
rect 1762 33182 1764 33234
rect 1708 33180 1764 33182
rect 1708 32508 1764 32564
rect 2828 40236 2884 40292
rect 3052 39506 3108 39508
rect 3052 39454 3054 39506
rect 3054 39454 3106 39506
rect 3106 39454 3108 39506
rect 3052 39452 3108 39454
rect 2940 38332 2996 38388
rect 2604 37490 2660 37492
rect 2604 37438 2606 37490
rect 2606 37438 2658 37490
rect 2658 37438 2660 37490
rect 2604 37436 2660 37438
rect 2828 37490 2884 37492
rect 2828 37438 2830 37490
rect 2830 37438 2882 37490
rect 2882 37438 2884 37490
rect 2828 37436 2884 37438
rect 2380 36316 2436 36372
rect 2716 36482 2772 36484
rect 2716 36430 2718 36482
rect 2718 36430 2770 36482
rect 2770 36430 2772 36482
rect 2716 36428 2772 36430
rect 3388 40236 3444 40292
rect 3612 40236 3668 40292
rect 4476 44714 4532 44716
rect 4476 44662 4478 44714
rect 4478 44662 4530 44714
rect 4530 44662 4532 44714
rect 4476 44660 4532 44662
rect 4580 44714 4636 44716
rect 4580 44662 4582 44714
rect 4582 44662 4634 44714
rect 4634 44662 4636 44714
rect 4580 44660 4636 44662
rect 4684 44714 4740 44716
rect 4684 44662 4686 44714
rect 4686 44662 4738 44714
rect 4738 44662 4740 44714
rect 4684 44660 4740 44662
rect 4844 43596 4900 43652
rect 5292 43650 5348 43652
rect 5292 43598 5294 43650
rect 5294 43598 5346 43650
rect 5346 43598 5348 43650
rect 5292 43596 5348 43598
rect 4060 43426 4116 43428
rect 4060 43374 4062 43426
rect 4062 43374 4114 43426
rect 4114 43374 4116 43426
rect 4060 43372 4116 43374
rect 4508 43260 4564 43316
rect 4476 43146 4532 43148
rect 4476 43094 4478 43146
rect 4478 43094 4530 43146
rect 4530 43094 4532 43146
rect 4476 43092 4532 43094
rect 4580 43146 4636 43148
rect 4580 43094 4582 43146
rect 4582 43094 4634 43146
rect 4634 43094 4636 43146
rect 4580 43092 4636 43094
rect 4684 43146 4740 43148
rect 4684 43094 4686 43146
rect 4686 43094 4738 43146
rect 4738 43094 4740 43146
rect 4684 43092 4740 43094
rect 5852 42252 5908 42308
rect 4060 41858 4116 41860
rect 4060 41806 4062 41858
rect 4062 41806 4114 41858
rect 4114 41806 4116 41858
rect 4060 41804 4116 41806
rect 4476 41578 4532 41580
rect 4476 41526 4478 41578
rect 4478 41526 4530 41578
rect 4530 41526 4532 41578
rect 4476 41524 4532 41526
rect 4580 41578 4636 41580
rect 4580 41526 4582 41578
rect 4582 41526 4634 41578
rect 4634 41526 4636 41578
rect 4580 41524 4636 41526
rect 4684 41578 4740 41580
rect 4684 41526 4686 41578
rect 4686 41526 4738 41578
rect 4738 41526 4740 41578
rect 4684 41524 4740 41526
rect 3948 39618 4004 39620
rect 3948 39566 3950 39618
rect 3950 39566 4002 39618
rect 4002 39566 4004 39618
rect 3948 39564 4004 39566
rect 4060 41132 4116 41188
rect 3500 39394 3556 39396
rect 3500 39342 3502 39394
rect 3502 39342 3554 39394
rect 3554 39342 3556 39394
rect 3500 39340 3556 39342
rect 3388 39228 3444 39284
rect 3612 39004 3668 39060
rect 3500 38946 3556 38948
rect 3500 38894 3502 38946
rect 3502 38894 3554 38946
rect 3554 38894 3556 38946
rect 3500 38892 3556 38894
rect 3836 38834 3892 38836
rect 3836 38782 3838 38834
rect 3838 38782 3890 38834
rect 3890 38782 3892 38834
rect 3836 38780 3892 38782
rect 3612 37548 3668 37604
rect 3836 38332 3892 38388
rect 3164 37154 3220 37156
rect 3164 37102 3166 37154
rect 3166 37102 3218 37154
rect 3218 37102 3220 37154
rect 3164 37100 3220 37102
rect 3164 36540 3220 36596
rect 3276 36482 3332 36484
rect 3276 36430 3278 36482
rect 3278 36430 3330 36482
rect 3330 36430 3332 36482
rect 3276 36428 3332 36430
rect 2828 36092 2884 36148
rect 2716 35756 2772 35812
rect 2604 35698 2660 35700
rect 2604 35646 2606 35698
rect 2606 35646 2658 35698
rect 2658 35646 2660 35698
rect 2604 35644 2660 35646
rect 2156 34860 2212 34916
rect 2044 34242 2100 34244
rect 2044 34190 2046 34242
rect 2046 34190 2098 34242
rect 2098 34190 2100 34242
rect 2044 34188 2100 34190
rect 2044 33122 2100 33124
rect 2044 33070 2046 33122
rect 2046 33070 2098 33122
rect 2098 33070 2100 33122
rect 2044 33068 2100 33070
rect 2044 31164 2100 31220
rect 1708 30716 1764 30772
rect 1484 28252 1540 28308
rect 1820 28364 1876 28420
rect 1708 27692 1764 27748
rect 1708 27132 1764 27188
rect 1708 25394 1764 25396
rect 1708 25342 1710 25394
rect 1710 25342 1762 25394
rect 1762 25342 1764 25394
rect 1708 25340 1764 25342
rect 1484 25004 1540 25060
rect 1708 23548 1764 23604
rect 1708 21756 1764 21812
rect 1708 19964 1764 20020
rect 1708 18172 1764 18228
rect 1708 16380 1764 16436
rect 2044 30098 2100 30100
rect 2044 30046 2046 30098
rect 2046 30046 2098 30098
rect 2098 30046 2100 30098
rect 2044 30044 2100 30046
rect 2044 28476 2100 28532
rect 3052 35532 3108 35588
rect 2604 34860 2660 34916
rect 2268 33292 2324 33348
rect 2492 33180 2548 33236
rect 2940 34636 2996 34692
rect 2828 34524 2884 34580
rect 3612 37212 3668 37268
rect 3948 38162 4004 38164
rect 3948 38110 3950 38162
rect 3950 38110 4002 38162
rect 4002 38110 4004 38162
rect 3948 38108 4004 38110
rect 4956 40460 5012 40516
rect 4476 40010 4532 40012
rect 4476 39958 4478 40010
rect 4478 39958 4530 40010
rect 4530 39958 4532 40010
rect 4476 39956 4532 39958
rect 4580 40010 4636 40012
rect 4580 39958 4582 40010
rect 4582 39958 4634 40010
rect 4634 39958 4636 40010
rect 4580 39956 4636 39958
rect 4684 40010 4740 40012
rect 4684 39958 4686 40010
rect 4686 39958 4738 40010
rect 4738 39958 4740 40010
rect 4684 39956 4740 39958
rect 5068 40348 5124 40404
rect 5740 40402 5796 40404
rect 5740 40350 5742 40402
rect 5742 40350 5794 40402
rect 5794 40350 5796 40402
rect 5740 40348 5796 40350
rect 4284 38834 4340 38836
rect 4284 38782 4286 38834
rect 4286 38782 4338 38834
rect 4338 38782 4340 38834
rect 4284 38780 4340 38782
rect 4476 38442 4532 38444
rect 4476 38390 4478 38442
rect 4478 38390 4530 38442
rect 4530 38390 4532 38442
rect 4476 38388 4532 38390
rect 4580 38442 4636 38444
rect 4580 38390 4582 38442
rect 4582 38390 4634 38442
rect 4634 38390 4636 38442
rect 4580 38388 4636 38390
rect 4684 38442 4740 38444
rect 4684 38390 4686 38442
rect 4686 38390 4738 38442
rect 4738 38390 4740 38442
rect 4684 38388 4740 38390
rect 4956 38274 5012 38276
rect 4956 38222 4958 38274
rect 4958 38222 5010 38274
rect 5010 38222 5012 38274
rect 4956 38220 5012 38222
rect 4732 38050 4788 38052
rect 4732 37998 4734 38050
rect 4734 37998 4786 38050
rect 4786 37998 4788 38050
rect 4732 37996 4788 37998
rect 3500 35586 3556 35588
rect 3500 35534 3502 35586
rect 3502 35534 3554 35586
rect 3554 35534 3556 35586
rect 3500 35532 3556 35534
rect 3948 37548 4004 37604
rect 4476 36874 4532 36876
rect 4476 36822 4478 36874
rect 4478 36822 4530 36874
rect 4530 36822 4532 36874
rect 4476 36820 4532 36822
rect 4580 36874 4636 36876
rect 4580 36822 4582 36874
rect 4582 36822 4634 36874
rect 4634 36822 4636 36874
rect 4580 36820 4636 36822
rect 4684 36874 4740 36876
rect 4684 36822 4686 36874
rect 4686 36822 4738 36874
rect 4738 36822 4740 36874
rect 4684 36820 4740 36822
rect 3164 34636 3220 34692
rect 3052 33516 3108 33572
rect 2828 33292 2884 33348
rect 2380 29932 2436 29988
rect 2380 28924 2436 28980
rect 2380 28642 2436 28644
rect 2380 28590 2382 28642
rect 2382 28590 2434 28642
rect 2434 28590 2436 28642
rect 2380 28588 2436 28590
rect 3164 33234 3220 33236
rect 3164 33182 3166 33234
rect 3166 33182 3218 33234
rect 3218 33182 3220 33234
rect 3164 33180 3220 33182
rect 2828 29260 2884 29316
rect 2940 31890 2996 31892
rect 2940 31838 2942 31890
rect 2942 31838 2994 31890
rect 2994 31838 2996 31890
rect 2940 31836 2996 31838
rect 3388 31724 3444 31780
rect 3052 31106 3108 31108
rect 3052 31054 3054 31106
rect 3054 31054 3106 31106
rect 3106 31054 3108 31106
rect 3052 31052 3108 31054
rect 3612 33122 3668 33124
rect 3612 33070 3614 33122
rect 3614 33070 3666 33122
rect 3666 33070 3668 33122
rect 3612 33068 3668 33070
rect 3948 35420 4004 35476
rect 4284 35980 4340 36036
rect 4620 35922 4676 35924
rect 4620 35870 4622 35922
rect 4622 35870 4674 35922
rect 4674 35870 4676 35922
rect 4620 35868 4676 35870
rect 4284 35532 4340 35588
rect 4476 35306 4532 35308
rect 4476 35254 4478 35306
rect 4478 35254 4530 35306
rect 4530 35254 4532 35306
rect 4476 35252 4532 35254
rect 4580 35306 4636 35308
rect 4580 35254 4582 35306
rect 4582 35254 4634 35306
rect 4634 35254 4636 35306
rect 4580 35252 4636 35254
rect 4684 35306 4740 35308
rect 4684 35254 4686 35306
rect 4686 35254 4738 35306
rect 4738 35254 4740 35306
rect 4844 35308 4900 35364
rect 4684 35252 4740 35254
rect 4396 34300 4452 34356
rect 4476 33738 4532 33740
rect 4476 33686 4478 33738
rect 4478 33686 4530 33738
rect 4530 33686 4532 33738
rect 4476 33684 4532 33686
rect 4580 33738 4636 33740
rect 4580 33686 4582 33738
rect 4582 33686 4634 33738
rect 4634 33686 4636 33738
rect 4580 33684 4636 33686
rect 4684 33738 4740 33740
rect 4684 33686 4686 33738
rect 4686 33686 4738 33738
rect 4738 33686 4740 33738
rect 4684 33684 4740 33686
rect 4620 33516 4676 33572
rect 5068 33346 5124 33348
rect 5068 33294 5070 33346
rect 5070 33294 5122 33346
rect 5122 33294 5124 33346
rect 5068 33292 5124 33294
rect 3724 32060 3780 32116
rect 4284 33180 4340 33236
rect 3612 31836 3668 31892
rect 3724 31724 3780 31780
rect 2940 28588 2996 28644
rect 2492 28418 2548 28420
rect 2492 28366 2494 28418
rect 2494 28366 2546 28418
rect 2546 28366 2548 28418
rect 2492 28364 2548 28366
rect 2716 28418 2772 28420
rect 2716 28366 2718 28418
rect 2718 28366 2770 28418
rect 2770 28366 2772 28418
rect 2716 28364 2772 28366
rect 2492 27746 2548 27748
rect 2492 27694 2494 27746
rect 2494 27694 2546 27746
rect 2546 27694 2548 27746
rect 2492 27692 2548 27694
rect 3164 29986 3220 29988
rect 3164 29934 3166 29986
rect 3166 29934 3218 29986
rect 3218 29934 3220 29986
rect 3164 29932 3220 29934
rect 3388 30882 3444 30884
rect 3388 30830 3390 30882
rect 3390 30830 3442 30882
rect 3442 30830 3444 30882
rect 3388 30828 3444 30830
rect 4060 32060 4116 32116
rect 3724 29820 3780 29876
rect 3164 29260 3220 29316
rect 2492 25394 2548 25396
rect 2492 25342 2494 25394
rect 2494 25342 2546 25394
rect 2546 25342 2548 25394
rect 2492 25340 2548 25342
rect 2044 23826 2100 23828
rect 2044 23774 2046 23826
rect 2046 23774 2098 23826
rect 2098 23774 2100 23826
rect 2044 23772 2100 23774
rect 3276 28530 3332 28532
rect 3276 28478 3278 28530
rect 3278 28478 3330 28530
rect 3330 28478 3332 28530
rect 3276 28476 3332 28478
rect 3948 28642 4004 28644
rect 3948 28590 3950 28642
rect 3950 28590 4002 28642
rect 4002 28590 4004 28642
rect 3948 28588 4004 28590
rect 3500 28418 3556 28420
rect 3500 28366 3502 28418
rect 3502 28366 3554 28418
rect 3554 28366 3556 28418
rect 3500 28364 3556 28366
rect 3388 26908 3444 26964
rect 3164 23772 3220 23828
rect 2492 23548 2548 23604
rect 2380 23436 2436 23492
rect 2492 21756 2548 21812
rect 2492 19964 2548 20020
rect 2492 18172 2548 18228
rect 2492 16380 2548 16436
rect 1820 15148 1876 15204
rect 1708 14588 1764 14644
rect 1708 12850 1764 12852
rect 1708 12798 1710 12850
rect 1710 12798 1762 12850
rect 1762 12798 1764 12850
rect 1708 12796 1764 12798
rect 1708 11004 1764 11060
rect 2492 14588 2548 14644
rect 2044 13356 2100 13412
rect 3948 28082 4004 28084
rect 3948 28030 3950 28082
rect 3950 28030 4002 28082
rect 4002 28030 4004 28082
rect 3948 28028 4004 28030
rect 5628 40236 5684 40292
rect 5292 39564 5348 39620
rect 5740 39452 5796 39508
rect 5852 39058 5908 39060
rect 5852 39006 5854 39058
rect 5854 39006 5906 39058
rect 5906 39006 5908 39058
rect 5852 39004 5908 39006
rect 5740 38946 5796 38948
rect 5740 38894 5742 38946
rect 5742 38894 5794 38946
rect 5794 38894 5796 38946
rect 5740 38892 5796 38894
rect 7420 48860 7476 48916
rect 6636 48300 6692 48356
rect 6412 47516 6468 47572
rect 7084 48354 7140 48356
rect 7084 48302 7086 48354
rect 7086 48302 7138 48354
rect 7138 48302 7140 48354
rect 7084 48300 7140 48302
rect 6188 45500 6244 45556
rect 6524 45388 6580 45444
rect 7308 47068 7364 47124
rect 7532 46620 7588 46676
rect 6748 45388 6804 45444
rect 7084 45612 7140 45668
rect 6188 40514 6244 40516
rect 6188 40462 6190 40514
rect 6190 40462 6242 40514
rect 6242 40462 6244 40514
rect 6188 40460 6244 40462
rect 6076 38892 6132 38948
rect 6972 45500 7028 45556
rect 6860 44156 6916 44212
rect 6860 43708 6916 43764
rect 6524 43650 6580 43652
rect 6524 43598 6526 43650
rect 6526 43598 6578 43650
rect 6578 43598 6580 43650
rect 6524 43596 6580 43598
rect 6636 42252 6692 42308
rect 6412 42082 6468 42084
rect 6412 42030 6414 42082
rect 6414 42030 6466 42082
rect 6466 42030 6468 42082
rect 6412 42028 6468 42030
rect 6412 39564 6468 39620
rect 6412 38668 6468 38724
rect 5628 37772 5684 37828
rect 5628 36316 5684 36372
rect 5404 35532 5460 35588
rect 5180 33180 5236 33236
rect 5292 34636 5348 34692
rect 5404 34354 5460 34356
rect 5404 34302 5406 34354
rect 5406 34302 5458 34354
rect 5458 34302 5460 34354
rect 5404 34300 5460 34302
rect 4956 32562 5012 32564
rect 4956 32510 4958 32562
rect 4958 32510 5010 32562
rect 5010 32510 5012 32562
rect 4956 32508 5012 32510
rect 4476 32170 4532 32172
rect 4476 32118 4478 32170
rect 4478 32118 4530 32170
rect 4530 32118 4532 32170
rect 4476 32116 4532 32118
rect 4580 32170 4636 32172
rect 4580 32118 4582 32170
rect 4582 32118 4634 32170
rect 4634 32118 4636 32170
rect 4580 32116 4636 32118
rect 4684 32170 4740 32172
rect 4684 32118 4686 32170
rect 4686 32118 4738 32170
rect 4738 32118 4740 32170
rect 4684 32116 4740 32118
rect 6748 41804 6804 41860
rect 6748 40348 6804 40404
rect 6748 38834 6804 38836
rect 6748 38782 6750 38834
rect 6750 38782 6802 38834
rect 6802 38782 6804 38834
rect 6748 38780 6804 38782
rect 7308 43708 7364 43764
rect 11788 55186 11844 55188
rect 11788 55134 11790 55186
rect 11790 55134 11842 55186
rect 11842 55134 11844 55186
rect 11788 55132 11844 55134
rect 13580 55298 13636 55300
rect 13580 55246 13582 55298
rect 13582 55246 13634 55298
rect 13634 55246 13636 55298
rect 13580 55244 13636 55246
rect 12684 55020 12740 55076
rect 12796 53788 12852 53844
rect 9884 53058 9940 53060
rect 9884 53006 9886 53058
rect 9886 53006 9938 53058
rect 9938 53006 9940 53058
rect 9884 53004 9940 53006
rect 11564 53506 11620 53508
rect 11564 53454 11566 53506
rect 11566 53454 11618 53506
rect 11618 53454 11620 53506
rect 11564 53452 11620 53454
rect 10556 53058 10612 53060
rect 10556 53006 10558 53058
rect 10558 53006 10610 53058
rect 10610 53006 10612 53058
rect 10556 53004 10612 53006
rect 10220 52556 10276 52612
rect 10444 52668 10500 52724
rect 10332 52444 10388 52500
rect 8988 51884 9044 51940
rect 10108 51772 10164 51828
rect 11116 53004 11172 53060
rect 10668 52946 10724 52948
rect 10668 52894 10670 52946
rect 10670 52894 10722 52946
rect 10722 52894 10724 52946
rect 10668 52892 10724 52894
rect 10892 52946 10948 52948
rect 10892 52894 10894 52946
rect 10894 52894 10946 52946
rect 10946 52894 10948 52946
rect 10892 52892 10948 52894
rect 11004 52722 11060 52724
rect 11004 52670 11006 52722
rect 11006 52670 11058 52722
rect 11058 52670 11060 52722
rect 11004 52668 11060 52670
rect 10780 51436 10836 51492
rect 10892 51548 10948 51604
rect 8988 51324 9044 51380
rect 12348 53116 12404 53172
rect 11340 52162 11396 52164
rect 11340 52110 11342 52162
rect 11342 52110 11394 52162
rect 11394 52110 11396 52162
rect 11340 52108 11396 52110
rect 11564 52892 11620 52948
rect 12796 53170 12852 53172
rect 12796 53118 12798 53170
rect 12798 53118 12850 53170
rect 12850 53118 12852 53170
rect 12796 53116 12852 53118
rect 13804 53116 13860 53172
rect 11676 52668 11732 52724
rect 12684 52556 12740 52612
rect 12348 52162 12404 52164
rect 12348 52110 12350 52162
rect 12350 52110 12402 52162
rect 12402 52110 12404 52162
rect 12348 52108 12404 52110
rect 11564 51436 11620 51492
rect 11116 49980 11172 50036
rect 10780 49868 10836 49924
rect 8204 48972 8260 49028
rect 8092 48860 8148 48916
rect 8988 49810 9044 49812
rect 8988 49758 8990 49810
rect 8990 49758 9042 49810
rect 9042 49758 9044 49810
rect 8988 49756 9044 49758
rect 12012 51602 12068 51604
rect 12012 51550 12014 51602
rect 12014 51550 12066 51602
rect 12066 51550 12068 51602
rect 12012 51548 12068 51550
rect 11900 51212 11956 51268
rect 12796 52444 12852 52500
rect 12012 50034 12068 50036
rect 12012 49982 12014 50034
rect 12014 49982 12066 50034
rect 12066 49982 12068 50034
rect 12012 49980 12068 49982
rect 12572 49980 12628 50036
rect 10556 49810 10612 49812
rect 10556 49758 10558 49810
rect 10558 49758 10610 49810
rect 10610 49758 10612 49810
rect 10556 49756 10612 49758
rect 8428 48860 8484 48916
rect 10108 49196 10164 49252
rect 8316 48412 8372 48468
rect 9660 48412 9716 48468
rect 8764 47458 8820 47460
rect 8764 47406 8766 47458
rect 8766 47406 8818 47458
rect 8818 47406 8820 47458
rect 8764 47404 8820 47406
rect 8316 47068 8372 47124
rect 8988 46844 9044 46900
rect 7868 46786 7924 46788
rect 7868 46734 7870 46786
rect 7870 46734 7922 46786
rect 7922 46734 7924 46786
rect 7868 46732 7924 46734
rect 7756 46620 7812 46676
rect 8092 45666 8148 45668
rect 8092 45614 8094 45666
rect 8094 45614 8146 45666
rect 8146 45614 8148 45666
rect 8092 45612 8148 45614
rect 7980 45388 8036 45444
rect 8652 45890 8708 45892
rect 8652 45838 8654 45890
rect 8654 45838 8706 45890
rect 8706 45838 8708 45890
rect 8652 45836 8708 45838
rect 8764 45724 8820 45780
rect 8316 45612 8372 45668
rect 7756 45106 7812 45108
rect 7756 45054 7758 45106
rect 7758 45054 7810 45106
rect 7810 45054 7812 45106
rect 7756 45052 7812 45054
rect 7980 44268 8036 44324
rect 8092 44210 8148 44212
rect 8092 44158 8094 44210
rect 8094 44158 8146 44210
rect 8146 44158 8148 44210
rect 8092 44156 8148 44158
rect 7980 43708 8036 43764
rect 7756 43650 7812 43652
rect 7756 43598 7758 43650
rect 7758 43598 7810 43650
rect 7810 43598 7812 43650
rect 7756 43596 7812 43598
rect 7868 43372 7924 43428
rect 7196 42028 7252 42084
rect 7868 42754 7924 42756
rect 7868 42702 7870 42754
rect 7870 42702 7922 42754
rect 7922 42702 7924 42754
rect 7868 42700 7924 42702
rect 7196 40460 7252 40516
rect 7644 42028 7700 42084
rect 8540 43708 8596 43764
rect 8316 42812 8372 42868
rect 8204 42588 8260 42644
rect 8092 40402 8148 40404
rect 8092 40350 8094 40402
rect 8094 40350 8146 40402
rect 8146 40350 8148 40402
rect 8092 40348 8148 40350
rect 8204 40236 8260 40292
rect 7756 39788 7812 39844
rect 7308 39564 7364 39620
rect 7420 39004 7476 39060
rect 5964 36370 6020 36372
rect 5964 36318 5966 36370
rect 5966 36318 6018 36370
rect 6018 36318 6020 36370
rect 5964 36316 6020 36318
rect 5740 35308 5796 35364
rect 5628 31948 5684 32004
rect 5516 31164 5572 31220
rect 4396 30828 4452 30884
rect 4476 30602 4532 30604
rect 4476 30550 4478 30602
rect 4478 30550 4530 30602
rect 4530 30550 4532 30602
rect 4476 30548 4532 30550
rect 4580 30602 4636 30604
rect 4580 30550 4582 30602
rect 4582 30550 4634 30602
rect 4634 30550 4636 30602
rect 4580 30548 4636 30550
rect 4684 30602 4740 30604
rect 4684 30550 4686 30602
rect 4686 30550 4738 30602
rect 4738 30550 4740 30602
rect 4684 30548 4740 30550
rect 5516 30994 5572 30996
rect 5516 30942 5518 30994
rect 5518 30942 5570 30994
rect 5570 30942 5572 30994
rect 5516 30940 5572 30942
rect 4172 29986 4228 29988
rect 4172 29934 4174 29986
rect 4174 29934 4226 29986
rect 4226 29934 4228 29986
rect 4172 29932 4228 29934
rect 4620 29426 4676 29428
rect 4620 29374 4622 29426
rect 4622 29374 4674 29426
rect 4674 29374 4676 29426
rect 4620 29372 4676 29374
rect 4476 29034 4532 29036
rect 4476 28982 4478 29034
rect 4478 28982 4530 29034
rect 4530 28982 4532 29034
rect 4476 28980 4532 28982
rect 4580 29034 4636 29036
rect 4580 28982 4582 29034
rect 4582 28982 4634 29034
rect 4634 28982 4636 29034
rect 4580 28980 4636 28982
rect 4684 29034 4740 29036
rect 4684 28982 4686 29034
rect 4686 28982 4738 29034
rect 4738 28982 4740 29034
rect 4684 28980 4740 28982
rect 4844 28252 4900 28308
rect 5068 29932 5124 29988
rect 6748 36370 6804 36372
rect 6748 36318 6750 36370
rect 6750 36318 6802 36370
rect 6802 36318 6804 36370
rect 6748 36316 6804 36318
rect 6300 35084 6356 35140
rect 6188 34690 6244 34692
rect 6188 34638 6190 34690
rect 6190 34638 6242 34690
rect 6242 34638 6244 34690
rect 6188 34636 6244 34638
rect 6636 34354 6692 34356
rect 6636 34302 6638 34354
rect 6638 34302 6690 34354
rect 6690 34302 6692 34354
rect 6636 34300 6692 34302
rect 6524 34188 6580 34244
rect 5964 33346 6020 33348
rect 5964 33294 5966 33346
rect 5966 33294 6018 33346
rect 6018 33294 6020 33346
rect 5964 33292 6020 33294
rect 6636 33516 6692 33572
rect 6636 32284 6692 32340
rect 6076 31276 6132 31332
rect 5964 30940 6020 30996
rect 5852 29986 5908 29988
rect 5852 29934 5854 29986
rect 5854 29934 5906 29986
rect 5906 29934 5908 29986
rect 5852 29932 5908 29934
rect 5628 29484 5684 29540
rect 6188 30098 6244 30100
rect 6188 30046 6190 30098
rect 6190 30046 6242 30098
rect 6242 30046 6244 30098
rect 6188 30044 6244 30046
rect 5068 29260 5124 29316
rect 5740 28588 5796 28644
rect 5292 28476 5348 28532
rect 5964 28364 6020 28420
rect 5292 28082 5348 28084
rect 5292 28030 5294 28082
rect 5294 28030 5346 28082
rect 5346 28030 5348 28082
rect 5292 28028 5348 28030
rect 4956 27916 5012 27972
rect 4284 27580 4340 27636
rect 4476 27466 4532 27468
rect 4476 27414 4478 27466
rect 4478 27414 4530 27466
rect 4530 27414 4532 27466
rect 4476 27412 4532 27414
rect 4580 27466 4636 27468
rect 4580 27414 4582 27466
rect 4582 27414 4634 27466
rect 4634 27414 4636 27466
rect 4580 27412 4636 27414
rect 4684 27466 4740 27468
rect 4684 27414 4686 27466
rect 4686 27414 4738 27466
rect 4738 27414 4740 27466
rect 4684 27412 4740 27414
rect 4476 25898 4532 25900
rect 4476 25846 4478 25898
rect 4478 25846 4530 25898
rect 4530 25846 4532 25898
rect 4476 25844 4532 25846
rect 4580 25898 4636 25900
rect 4580 25846 4582 25898
rect 4582 25846 4634 25898
rect 4634 25846 4636 25898
rect 4580 25844 4636 25846
rect 4684 25898 4740 25900
rect 4684 25846 4686 25898
rect 4686 25846 4738 25898
rect 4738 25846 4740 25898
rect 4684 25844 4740 25846
rect 5852 28252 5908 28308
rect 5404 27804 5460 27860
rect 5516 27692 5572 27748
rect 6636 30098 6692 30100
rect 6636 30046 6638 30098
rect 6638 30046 6690 30098
rect 6690 30046 6692 30098
rect 6636 30044 6692 30046
rect 6412 29820 6468 29876
rect 5964 27692 6020 27748
rect 5964 27074 6020 27076
rect 5964 27022 5966 27074
rect 5966 27022 6018 27074
rect 6018 27022 6020 27074
rect 5964 27020 6020 27022
rect 5740 26908 5796 26964
rect 4732 25004 4788 25060
rect 4476 24330 4532 24332
rect 4476 24278 4478 24330
rect 4478 24278 4530 24330
rect 4530 24278 4532 24330
rect 4476 24276 4532 24278
rect 4580 24330 4636 24332
rect 4580 24278 4582 24330
rect 4582 24278 4634 24330
rect 4634 24278 4636 24330
rect 4580 24276 4636 24278
rect 4684 24330 4740 24332
rect 4684 24278 4686 24330
rect 4686 24278 4738 24330
rect 4738 24278 4740 24330
rect 4684 24276 4740 24278
rect 6412 27916 6468 27972
rect 6076 26460 6132 26516
rect 5964 26290 6020 26292
rect 5964 26238 5966 26290
rect 5966 26238 6018 26290
rect 6018 26238 6020 26290
rect 5964 26236 6020 26238
rect 5852 23212 5908 23268
rect 4476 22762 4532 22764
rect 4476 22710 4478 22762
rect 4478 22710 4530 22762
rect 4530 22710 4532 22762
rect 4476 22708 4532 22710
rect 4580 22762 4636 22764
rect 4580 22710 4582 22762
rect 4582 22710 4634 22762
rect 4634 22710 4636 22762
rect 4580 22708 4636 22710
rect 4684 22762 4740 22764
rect 4684 22710 4686 22762
rect 4686 22710 4738 22762
rect 4738 22710 4740 22762
rect 4684 22708 4740 22710
rect 4476 21194 4532 21196
rect 4476 21142 4478 21194
rect 4478 21142 4530 21194
rect 4530 21142 4532 21194
rect 4476 21140 4532 21142
rect 4580 21194 4636 21196
rect 4580 21142 4582 21194
rect 4582 21142 4634 21194
rect 4634 21142 4636 21194
rect 4580 21140 4636 21142
rect 4684 21194 4740 21196
rect 4684 21142 4686 21194
rect 4686 21142 4738 21194
rect 4738 21142 4740 21194
rect 4684 21140 4740 21142
rect 4476 19626 4532 19628
rect 4476 19574 4478 19626
rect 4478 19574 4530 19626
rect 4530 19574 4532 19626
rect 4476 19572 4532 19574
rect 4580 19626 4636 19628
rect 4580 19574 4582 19626
rect 4582 19574 4634 19626
rect 4634 19574 4636 19626
rect 4580 19572 4636 19574
rect 4684 19626 4740 19628
rect 4684 19574 4686 19626
rect 4686 19574 4738 19626
rect 4738 19574 4740 19626
rect 4684 19572 4740 19574
rect 4476 18058 4532 18060
rect 4476 18006 4478 18058
rect 4478 18006 4530 18058
rect 4530 18006 4532 18058
rect 4476 18004 4532 18006
rect 4580 18058 4636 18060
rect 4580 18006 4582 18058
rect 4582 18006 4634 18058
rect 4634 18006 4636 18058
rect 4580 18004 4636 18006
rect 4684 18058 4740 18060
rect 4684 18006 4686 18058
rect 4686 18006 4738 18058
rect 4738 18006 4740 18058
rect 4684 18004 4740 18006
rect 4476 16490 4532 16492
rect 4476 16438 4478 16490
rect 4478 16438 4530 16490
rect 4530 16438 4532 16490
rect 4476 16436 4532 16438
rect 4580 16490 4636 16492
rect 4580 16438 4582 16490
rect 4582 16438 4634 16490
rect 4634 16438 4636 16490
rect 4580 16436 4636 16438
rect 4684 16490 4740 16492
rect 4684 16438 4686 16490
rect 4686 16438 4738 16490
rect 4738 16438 4740 16490
rect 4684 16436 4740 16438
rect 4476 14922 4532 14924
rect 4476 14870 4478 14922
rect 4478 14870 4530 14922
rect 4530 14870 4532 14922
rect 4476 14868 4532 14870
rect 4580 14922 4636 14924
rect 4580 14870 4582 14922
rect 4582 14870 4634 14922
rect 4634 14870 4636 14922
rect 4580 14868 4636 14870
rect 4684 14922 4740 14924
rect 4684 14870 4686 14922
rect 4686 14870 4738 14922
rect 4738 14870 4740 14922
rect 4684 14868 4740 14870
rect 3836 13356 3892 13412
rect 4476 13354 4532 13356
rect 4476 13302 4478 13354
rect 4478 13302 4530 13354
rect 4530 13302 4532 13354
rect 4476 13300 4532 13302
rect 4580 13354 4636 13356
rect 4580 13302 4582 13354
rect 4582 13302 4634 13354
rect 4634 13302 4636 13354
rect 4580 13300 4636 13302
rect 4684 13354 4740 13356
rect 4684 13302 4686 13354
rect 4686 13302 4738 13354
rect 4738 13302 4740 13354
rect 4684 13300 4740 13302
rect 2492 12850 2548 12852
rect 2492 12798 2494 12850
rect 2494 12798 2546 12850
rect 2546 12798 2548 12850
rect 2492 12796 2548 12798
rect 4476 11786 4532 11788
rect 4476 11734 4478 11786
rect 4478 11734 4530 11786
rect 4530 11734 4532 11786
rect 4476 11732 4532 11734
rect 4580 11786 4636 11788
rect 4580 11734 4582 11786
rect 4582 11734 4634 11786
rect 4634 11734 4636 11786
rect 4580 11732 4636 11734
rect 4684 11786 4740 11788
rect 4684 11734 4686 11786
rect 4686 11734 4738 11786
rect 4738 11734 4740 11786
rect 4684 11732 4740 11734
rect 2044 11282 2100 11284
rect 2044 11230 2046 11282
rect 2046 11230 2098 11282
rect 2098 11230 2100 11282
rect 2044 11228 2100 11230
rect 6300 11228 6356 11284
rect 2492 11004 2548 11060
rect 4476 10218 4532 10220
rect 4476 10166 4478 10218
rect 4478 10166 4530 10218
rect 4530 10166 4532 10218
rect 4476 10164 4532 10166
rect 4580 10218 4636 10220
rect 4580 10166 4582 10218
rect 4582 10166 4634 10218
rect 4634 10166 4636 10218
rect 4580 10164 4636 10166
rect 4684 10218 4740 10220
rect 4684 10166 4686 10218
rect 4686 10166 4738 10218
rect 4738 10166 4740 10218
rect 4684 10164 4740 10166
rect 2380 9996 2436 10052
rect 1708 9212 1764 9268
rect 1708 7980 1764 8036
rect 1708 7420 1764 7476
rect 1260 5852 1316 5908
rect 2156 5852 2212 5908
rect 1708 5628 1764 5684
rect 2044 4562 2100 4564
rect 2044 4510 2046 4562
rect 2046 4510 2098 4562
rect 2098 4510 2100 4562
rect 2044 4508 2100 4510
rect 1708 3836 1764 3892
rect 6748 27132 6804 27188
rect 6860 25676 6916 25732
rect 7756 39004 7812 39060
rect 8092 40124 8148 40180
rect 8764 42754 8820 42756
rect 8764 42702 8766 42754
rect 8766 42702 8818 42754
rect 8818 42702 8820 42754
rect 8764 42700 8820 42702
rect 9100 46732 9156 46788
rect 9884 46002 9940 46004
rect 9884 45950 9886 46002
rect 9886 45950 9938 46002
rect 9938 45950 9940 46002
rect 9884 45948 9940 45950
rect 9548 45836 9604 45892
rect 9324 45778 9380 45780
rect 9324 45726 9326 45778
rect 9326 45726 9378 45778
rect 9378 45726 9380 45778
rect 9324 45724 9380 45726
rect 8876 42642 8932 42644
rect 8876 42590 8878 42642
rect 8878 42590 8930 42642
rect 8930 42590 8932 42642
rect 8876 42588 8932 42590
rect 8876 42194 8932 42196
rect 8876 42142 8878 42194
rect 8878 42142 8930 42194
rect 8930 42142 8932 42194
rect 8876 42140 8932 42142
rect 9324 42700 9380 42756
rect 9436 41804 9492 41860
rect 8764 40460 8820 40516
rect 7084 37772 7140 37828
rect 7420 37154 7476 37156
rect 7420 37102 7422 37154
rect 7422 37102 7474 37154
rect 7474 37102 7476 37154
rect 7420 37100 7476 37102
rect 8204 39788 8260 39844
rect 7980 39618 8036 39620
rect 7980 39566 7982 39618
rect 7982 39566 8034 39618
rect 8034 39566 8036 39618
rect 7980 39564 8036 39566
rect 8316 39676 8372 39732
rect 8092 38722 8148 38724
rect 8092 38670 8094 38722
rect 8094 38670 8146 38722
rect 8146 38670 8148 38722
rect 8092 38668 8148 38670
rect 8204 37996 8260 38052
rect 8652 38722 8708 38724
rect 8652 38670 8654 38722
rect 8654 38670 8706 38722
rect 8706 38670 8708 38722
rect 8652 38668 8708 38670
rect 8988 37324 9044 37380
rect 8428 37100 8484 37156
rect 7756 36092 7812 36148
rect 7532 33964 7588 34020
rect 7084 33180 7140 33236
rect 7308 32562 7364 32564
rect 7308 32510 7310 32562
rect 7310 32510 7362 32562
rect 7362 32510 7364 32562
rect 7308 32508 7364 32510
rect 7084 31948 7140 32004
rect 8204 35308 8260 35364
rect 8988 36988 9044 37044
rect 8988 35756 9044 35812
rect 8540 35644 8596 35700
rect 7868 34636 7924 34692
rect 8092 34412 8148 34468
rect 7644 32956 7700 33012
rect 7420 31276 7476 31332
rect 7532 31218 7588 31220
rect 7532 31166 7534 31218
rect 7534 31166 7586 31218
rect 7586 31166 7588 31218
rect 7532 31164 7588 31166
rect 7980 30268 8036 30324
rect 7756 29986 7812 29988
rect 7756 29934 7758 29986
rect 7758 29934 7810 29986
rect 7810 29934 7812 29986
rect 7756 29932 7812 29934
rect 7868 29820 7924 29876
rect 7532 29708 7588 29764
rect 7420 29538 7476 29540
rect 7420 29486 7422 29538
rect 7422 29486 7474 29538
rect 7474 29486 7476 29538
rect 7420 29484 7476 29486
rect 7756 28476 7812 28532
rect 7084 27858 7140 27860
rect 7084 27806 7086 27858
rect 7086 27806 7138 27858
rect 7138 27806 7140 27858
rect 7084 27804 7140 27806
rect 7756 27858 7812 27860
rect 7756 27806 7758 27858
rect 7758 27806 7810 27858
rect 7810 27806 7812 27858
rect 7756 27804 7812 27806
rect 7980 27468 8036 27524
rect 7868 26402 7924 26404
rect 7868 26350 7870 26402
rect 7870 26350 7922 26402
rect 7922 26350 7924 26402
rect 7868 26348 7924 26350
rect 7644 26236 7700 26292
rect 7308 25730 7364 25732
rect 7308 25678 7310 25730
rect 7310 25678 7362 25730
rect 7362 25678 7364 25730
rect 7308 25676 7364 25678
rect 7084 25618 7140 25620
rect 7084 25566 7086 25618
rect 7086 25566 7138 25618
rect 7138 25566 7140 25618
rect 7084 25564 7140 25566
rect 7532 25506 7588 25508
rect 7532 25454 7534 25506
rect 7534 25454 7586 25506
rect 7586 25454 7588 25506
rect 7532 25452 7588 25454
rect 7756 25564 7812 25620
rect 7868 25228 7924 25284
rect 7980 21756 8036 21812
rect 8540 34300 8596 34356
rect 8204 33964 8260 34020
rect 8652 33292 8708 33348
rect 8876 32844 8932 32900
rect 10556 49532 10612 49588
rect 10220 48300 10276 48356
rect 10332 46844 10388 46900
rect 11228 49586 11284 49588
rect 11228 49534 11230 49586
rect 11230 49534 11282 49586
rect 11282 49534 11284 49586
rect 11228 49532 11284 49534
rect 11116 49250 11172 49252
rect 11116 49198 11118 49250
rect 11118 49198 11170 49250
rect 11170 49198 11172 49250
rect 11116 49196 11172 49198
rect 10668 48748 10724 48804
rect 11340 48748 11396 48804
rect 10556 48242 10612 48244
rect 10556 48190 10558 48242
rect 10558 48190 10610 48242
rect 10610 48190 10612 48242
rect 10556 48188 10612 48190
rect 11452 48300 11508 48356
rect 11340 47740 11396 47796
rect 10780 47458 10836 47460
rect 10780 47406 10782 47458
rect 10782 47406 10834 47458
rect 10834 47406 10836 47458
rect 10780 47404 10836 47406
rect 11004 45948 11060 46004
rect 10892 45836 10948 45892
rect 10444 45666 10500 45668
rect 10444 45614 10446 45666
rect 10446 45614 10498 45666
rect 10498 45614 10500 45666
rect 10444 45612 10500 45614
rect 10780 45612 10836 45668
rect 10444 44828 10500 44884
rect 10556 44716 10612 44772
rect 10444 44322 10500 44324
rect 10444 44270 10446 44322
rect 10446 44270 10498 44322
rect 10498 44270 10500 44322
rect 10444 44268 10500 44270
rect 9996 43932 10052 43988
rect 9548 41298 9604 41300
rect 9548 41246 9550 41298
rect 9550 41246 9602 41298
rect 9602 41246 9604 41298
rect 9548 41244 9604 41246
rect 10108 43538 10164 43540
rect 10108 43486 10110 43538
rect 10110 43486 10162 43538
rect 10162 43486 10164 43538
rect 10108 43484 10164 43486
rect 9996 43426 10052 43428
rect 9996 43374 9998 43426
rect 9998 43374 10050 43426
rect 10050 43374 10052 43426
rect 9996 43372 10052 43374
rect 9772 42700 9828 42756
rect 9660 42252 9716 42308
rect 9548 41020 9604 41076
rect 9884 41244 9940 41300
rect 9884 40460 9940 40516
rect 9212 38220 9268 38276
rect 9436 38556 9492 38612
rect 9212 37324 9268 37380
rect 9212 33404 9268 33460
rect 9100 31836 9156 31892
rect 8428 31612 8484 31668
rect 9100 31388 9156 31444
rect 8988 30940 9044 30996
rect 8652 30044 8708 30100
rect 8540 29260 8596 29316
rect 8652 28588 8708 28644
rect 8876 28588 8932 28644
rect 8540 28252 8596 28308
rect 8764 28364 8820 28420
rect 8652 28082 8708 28084
rect 8652 28030 8654 28082
rect 8654 28030 8706 28082
rect 8706 28030 8708 28082
rect 8652 28028 8708 28030
rect 8876 28252 8932 28308
rect 8540 27468 8596 27524
rect 8652 27692 8708 27748
rect 9772 38220 9828 38276
rect 10444 43036 10500 43092
rect 10556 43820 10612 43876
rect 10332 42530 10388 42532
rect 10332 42478 10334 42530
rect 10334 42478 10386 42530
rect 10386 42478 10388 42530
rect 10332 42476 10388 42478
rect 11676 48018 11732 48020
rect 11676 47966 11678 48018
rect 11678 47966 11730 48018
rect 11730 47966 11732 48018
rect 11676 47964 11732 47966
rect 11788 47516 11844 47572
rect 11452 46674 11508 46676
rect 11452 46622 11454 46674
rect 11454 46622 11506 46674
rect 11506 46622 11508 46674
rect 11452 46620 11508 46622
rect 11340 45724 11396 45780
rect 11116 44716 11172 44772
rect 11228 44828 11284 44884
rect 11004 44322 11060 44324
rect 11004 44270 11006 44322
rect 11006 44270 11058 44322
rect 11058 44270 11060 44322
rect 11004 44268 11060 44270
rect 11004 43650 11060 43652
rect 11004 43598 11006 43650
rect 11006 43598 11058 43650
rect 11058 43598 11060 43650
rect 11004 43596 11060 43598
rect 10780 42754 10836 42756
rect 10780 42702 10782 42754
rect 10782 42702 10834 42754
rect 10834 42702 10836 42754
rect 10780 42700 10836 42702
rect 10892 42588 10948 42644
rect 10332 39788 10388 39844
rect 10556 40684 10612 40740
rect 10556 40348 10612 40404
rect 10332 39564 10388 39620
rect 10556 39228 10612 39284
rect 11452 45612 11508 45668
rect 11340 43708 11396 43764
rect 11452 43314 11508 43316
rect 11452 43262 11454 43314
rect 11454 43262 11506 43314
rect 11506 43262 11508 43314
rect 11452 43260 11508 43262
rect 11340 43036 11396 43092
rect 11340 42364 11396 42420
rect 11452 40684 11508 40740
rect 11452 40402 11508 40404
rect 11452 40350 11454 40402
rect 11454 40350 11506 40402
rect 11506 40350 11508 40402
rect 11452 40348 11508 40350
rect 11676 43708 11732 43764
rect 12796 48860 12852 48916
rect 12460 48802 12516 48804
rect 12460 48750 12462 48802
rect 12462 48750 12514 48802
rect 12514 48750 12516 48802
rect 12460 48748 12516 48750
rect 12124 47516 12180 47572
rect 12908 48748 12964 48804
rect 12012 45948 12068 46004
rect 12572 46508 12628 46564
rect 12124 45724 12180 45780
rect 11788 43372 11844 43428
rect 12124 43596 12180 43652
rect 11900 43260 11956 43316
rect 11788 42588 11844 42644
rect 12460 43426 12516 43428
rect 12460 43374 12462 43426
rect 12462 43374 12514 43426
rect 12514 43374 12516 43426
rect 12460 43372 12516 43374
rect 12236 42252 12292 42308
rect 12236 40908 12292 40964
rect 11676 40514 11732 40516
rect 11676 40462 11678 40514
rect 11678 40462 11730 40514
rect 11730 40462 11732 40514
rect 11676 40460 11732 40462
rect 10780 39618 10836 39620
rect 10780 39566 10782 39618
rect 10782 39566 10834 39618
rect 10834 39566 10836 39618
rect 10780 39564 10836 39566
rect 10780 38780 10836 38836
rect 9660 36988 9716 37044
rect 9772 35420 9828 35476
rect 10108 37266 10164 37268
rect 10108 37214 10110 37266
rect 10110 37214 10162 37266
rect 10162 37214 10164 37266
rect 10108 37212 10164 37214
rect 10332 36204 10388 36260
rect 10108 35922 10164 35924
rect 10108 35870 10110 35922
rect 10110 35870 10162 35922
rect 10162 35870 10164 35922
rect 10108 35868 10164 35870
rect 10556 37996 10612 38052
rect 10668 37660 10724 37716
rect 10556 36258 10612 36260
rect 10556 36206 10558 36258
rect 10558 36206 10610 36258
rect 10610 36206 10612 36258
rect 10556 36204 10612 36206
rect 11004 39394 11060 39396
rect 11004 39342 11006 39394
rect 11006 39342 11058 39394
rect 11058 39342 11060 39394
rect 11004 39340 11060 39342
rect 11228 39116 11284 39172
rect 11228 38274 11284 38276
rect 11228 38222 11230 38274
rect 11230 38222 11282 38274
rect 11282 38222 11284 38274
rect 11228 38220 11284 38222
rect 11116 37660 11172 37716
rect 11116 36988 11172 37044
rect 11116 36204 11172 36260
rect 10444 35644 10500 35700
rect 9884 35026 9940 35028
rect 9884 34974 9886 35026
rect 9886 34974 9938 35026
rect 9938 34974 9940 35026
rect 9884 34972 9940 34974
rect 9660 34524 9716 34580
rect 9660 34300 9716 34356
rect 9660 33458 9716 33460
rect 9660 33406 9662 33458
rect 9662 33406 9714 33458
rect 9714 33406 9716 33458
rect 9660 33404 9716 33406
rect 9548 31836 9604 31892
rect 9660 32844 9716 32900
rect 9436 31388 9492 31444
rect 9100 28812 9156 28868
rect 8988 27692 9044 27748
rect 9212 27186 9268 27188
rect 9212 27134 9214 27186
rect 9214 27134 9266 27186
rect 9266 27134 9268 27186
rect 9212 27132 9268 27134
rect 9100 27074 9156 27076
rect 9100 27022 9102 27074
rect 9102 27022 9154 27074
rect 9154 27022 9156 27074
rect 9100 27020 9156 27022
rect 9324 26850 9380 26852
rect 9324 26798 9326 26850
rect 9326 26798 9378 26850
rect 9378 26798 9380 26850
rect 9324 26796 9380 26798
rect 9660 29820 9716 29876
rect 9660 29426 9716 29428
rect 9660 29374 9662 29426
rect 9662 29374 9714 29426
rect 9714 29374 9716 29426
rect 9660 29372 9716 29374
rect 9772 28028 9828 28084
rect 9772 26908 9828 26964
rect 9548 26796 9604 26852
rect 9660 26514 9716 26516
rect 9660 26462 9662 26514
rect 9662 26462 9714 26514
rect 9714 26462 9716 26514
rect 9660 26460 9716 26462
rect 10220 35252 10276 35308
rect 10108 34300 10164 34356
rect 10108 34018 10164 34020
rect 10108 33966 10110 34018
rect 10110 33966 10162 34018
rect 10162 33966 10164 34018
rect 10108 33964 10164 33966
rect 10108 32172 10164 32228
rect 10108 30994 10164 30996
rect 10108 30942 10110 30994
rect 10110 30942 10162 30994
rect 10162 30942 10164 30994
rect 10108 30940 10164 30942
rect 9996 29932 10052 29988
rect 10556 35420 10612 35476
rect 10780 35420 10836 35476
rect 10556 34242 10612 34244
rect 10556 34190 10558 34242
rect 10558 34190 10610 34242
rect 10610 34190 10612 34242
rect 10556 34188 10612 34190
rect 10668 33964 10724 34020
rect 10444 33404 10500 33460
rect 10780 33404 10836 33460
rect 10668 33068 10724 33124
rect 10444 32562 10500 32564
rect 10444 32510 10446 32562
rect 10446 32510 10498 32562
rect 10498 32510 10500 32562
rect 10444 32508 10500 32510
rect 10892 32620 10948 32676
rect 11116 34188 11172 34244
rect 11116 33740 11172 33796
rect 11004 32284 11060 32340
rect 10892 31612 10948 31668
rect 11004 31388 11060 31444
rect 11340 34636 11396 34692
rect 11788 40236 11844 40292
rect 12124 40796 12180 40852
rect 12684 43932 12740 43988
rect 12684 43708 12740 43764
rect 12796 46732 12852 46788
rect 16828 55298 16884 55300
rect 16828 55246 16830 55298
rect 16830 55246 16882 55298
rect 16882 55246 16884 55298
rect 16828 55244 16884 55246
rect 14588 52220 14644 52276
rect 14812 52444 14868 52500
rect 13244 51884 13300 51940
rect 15484 53004 15540 53060
rect 15372 52444 15428 52500
rect 16044 53788 16100 53844
rect 15596 51996 15652 52052
rect 15148 51884 15204 51940
rect 15708 51938 15764 51940
rect 15708 51886 15710 51938
rect 15710 51886 15762 51938
rect 15762 51886 15764 51938
rect 15708 51884 15764 51886
rect 15036 51548 15092 51604
rect 16156 52892 16212 52948
rect 16492 52668 16548 52724
rect 16156 52220 16212 52276
rect 16268 52162 16324 52164
rect 16268 52110 16270 52162
rect 16270 52110 16322 52162
rect 16322 52110 16324 52162
rect 16268 52108 16324 52110
rect 16492 52108 16548 52164
rect 18508 55356 18564 55412
rect 17724 55298 17780 55300
rect 17724 55246 17726 55298
rect 17726 55246 17778 55298
rect 17778 55246 17780 55298
rect 17724 55244 17780 55246
rect 17836 54514 17892 54516
rect 17836 54462 17838 54514
rect 17838 54462 17890 54514
rect 17890 54462 17892 54514
rect 17836 54460 17892 54462
rect 18172 53506 18228 53508
rect 18172 53454 18174 53506
rect 18174 53454 18226 53506
rect 18226 53454 18228 53506
rect 18172 53452 18228 53454
rect 17276 52892 17332 52948
rect 17388 51996 17444 52052
rect 15820 51100 15876 51156
rect 13244 50428 13300 50484
rect 15596 50540 15652 50596
rect 13132 50034 13188 50036
rect 13132 49982 13134 50034
rect 13134 49982 13186 50034
rect 13186 49982 13188 50034
rect 13132 49980 13188 49982
rect 15372 49026 15428 49028
rect 15372 48974 15374 49026
rect 15374 48974 15426 49026
rect 15426 48974 15428 49026
rect 15372 48972 15428 48974
rect 13356 47628 13412 47684
rect 13132 47404 13188 47460
rect 13356 46898 13412 46900
rect 13356 46846 13358 46898
rect 13358 46846 13410 46898
rect 13410 46846 13412 46898
rect 13356 46844 13412 46846
rect 13132 46786 13188 46788
rect 13132 46734 13134 46786
rect 13134 46734 13186 46786
rect 13186 46734 13188 46786
rect 13132 46732 13188 46734
rect 13580 47292 13636 47348
rect 13916 48018 13972 48020
rect 13916 47966 13918 48018
rect 13918 47966 13970 48018
rect 13970 47966 13972 48018
rect 13916 47964 13972 47966
rect 14028 47458 14084 47460
rect 14028 47406 14030 47458
rect 14030 47406 14082 47458
rect 14082 47406 14084 47458
rect 14028 47404 14084 47406
rect 14028 46620 14084 46676
rect 14252 47516 14308 47572
rect 14476 48076 14532 48132
rect 14476 47628 14532 47684
rect 14812 47458 14868 47460
rect 14812 47406 14814 47458
rect 14814 47406 14866 47458
rect 14866 47406 14868 47458
rect 14812 47404 14868 47406
rect 14700 47292 14756 47348
rect 14476 47068 14532 47124
rect 14476 46060 14532 46116
rect 15260 48130 15316 48132
rect 15260 48078 15262 48130
rect 15262 48078 15314 48130
rect 15314 48078 15316 48130
rect 15260 48076 15316 48078
rect 15372 47458 15428 47460
rect 15372 47406 15374 47458
rect 15374 47406 15426 47458
rect 15426 47406 15428 47458
rect 15372 47404 15428 47406
rect 15820 47964 15876 48020
rect 15484 47068 15540 47124
rect 15036 46674 15092 46676
rect 15036 46622 15038 46674
rect 15038 46622 15090 46674
rect 15090 46622 15092 46674
rect 15036 46620 15092 46622
rect 13020 44380 13076 44436
rect 12684 43036 12740 43092
rect 12236 39564 12292 39620
rect 12348 38834 12404 38836
rect 12348 38782 12350 38834
rect 12350 38782 12402 38834
rect 12402 38782 12404 38834
rect 12348 38780 12404 38782
rect 11900 37324 11956 37380
rect 12124 38220 12180 38276
rect 12236 38162 12292 38164
rect 12236 38110 12238 38162
rect 12238 38110 12290 38162
rect 12290 38110 12292 38162
rect 12236 38108 12292 38110
rect 12124 37826 12180 37828
rect 12124 37774 12126 37826
rect 12126 37774 12178 37826
rect 12178 37774 12180 37826
rect 12124 37772 12180 37774
rect 12348 37772 12404 37828
rect 13804 45106 13860 45108
rect 13804 45054 13806 45106
rect 13806 45054 13858 45106
rect 13858 45054 13860 45106
rect 13804 45052 13860 45054
rect 13132 43650 13188 43652
rect 13132 43598 13134 43650
rect 13134 43598 13186 43650
rect 13186 43598 13188 43650
rect 13132 43596 13188 43598
rect 14476 44492 14532 44548
rect 13916 43538 13972 43540
rect 13916 43486 13918 43538
rect 13918 43486 13970 43538
rect 13970 43486 13972 43538
rect 13916 43484 13972 43486
rect 13468 43260 13524 43316
rect 13020 41244 13076 41300
rect 12908 40290 12964 40292
rect 12908 40238 12910 40290
rect 12910 40238 12962 40290
rect 12962 40238 12964 40290
rect 12908 40236 12964 40238
rect 12796 39452 12852 39508
rect 13580 41074 13636 41076
rect 13580 41022 13582 41074
rect 13582 41022 13634 41074
rect 13634 41022 13636 41074
rect 13580 41020 13636 41022
rect 13356 40684 13412 40740
rect 13132 39228 13188 39284
rect 13020 39058 13076 39060
rect 13020 39006 13022 39058
rect 13022 39006 13074 39058
rect 13074 39006 13076 39058
rect 13020 39004 13076 39006
rect 13804 42252 13860 42308
rect 12796 38108 12852 38164
rect 13356 38444 13412 38500
rect 13020 37884 13076 37940
rect 12124 36988 12180 37044
rect 12012 36092 12068 36148
rect 12012 35922 12068 35924
rect 12012 35870 12014 35922
rect 12014 35870 12066 35922
rect 12066 35870 12068 35922
rect 12012 35868 12068 35870
rect 12012 35644 12068 35700
rect 11564 35084 11620 35140
rect 11564 34802 11620 34804
rect 11564 34750 11566 34802
rect 11566 34750 11618 34802
rect 11618 34750 11620 34802
rect 11564 34748 11620 34750
rect 12012 34412 12068 34468
rect 11676 34300 11732 34356
rect 12236 35084 12292 35140
rect 12908 37660 12964 37716
rect 13244 37660 13300 37716
rect 12572 37324 12628 37380
rect 12908 37212 12964 37268
rect 12908 36428 12964 36484
rect 12572 36204 12628 36260
rect 13132 36092 13188 36148
rect 12572 34914 12628 34916
rect 12572 34862 12574 34914
rect 12574 34862 12626 34914
rect 12626 34862 12628 34914
rect 12572 34860 12628 34862
rect 12012 34018 12068 34020
rect 12012 33966 12014 34018
rect 12014 33966 12066 34018
rect 12066 33966 12068 34018
rect 12012 33964 12068 33966
rect 11452 30492 11508 30548
rect 11228 30380 11284 30436
rect 11564 30380 11620 30436
rect 10444 29932 10500 29988
rect 10668 29820 10724 29876
rect 10892 29932 10948 29988
rect 10668 29372 10724 29428
rect 10556 28588 10612 28644
rect 10108 27804 10164 27860
rect 9996 27746 10052 27748
rect 9996 27694 9998 27746
rect 9998 27694 10050 27746
rect 10050 27694 10052 27746
rect 9996 27692 10052 27694
rect 10108 26962 10164 26964
rect 10108 26910 10110 26962
rect 10110 26910 10162 26962
rect 10162 26910 10164 26962
rect 10108 26908 10164 26910
rect 9884 26460 9940 26516
rect 10220 26348 10276 26404
rect 9548 25676 9604 25732
rect 9660 26236 9716 26292
rect 9660 25564 9716 25620
rect 10220 25506 10276 25508
rect 10220 25454 10222 25506
rect 10222 25454 10274 25506
rect 10274 25454 10276 25506
rect 10220 25452 10276 25454
rect 9548 25394 9604 25396
rect 9548 25342 9550 25394
rect 9550 25342 9602 25394
rect 9602 25342 9604 25394
rect 9548 25340 9604 25342
rect 8204 25004 8260 25060
rect 8316 25228 8372 25284
rect 9884 23996 9940 24052
rect 11004 29426 11060 29428
rect 11004 29374 11006 29426
rect 11006 29374 11058 29426
rect 11058 29374 11060 29426
rect 11004 29372 11060 29374
rect 10892 28418 10948 28420
rect 10892 28366 10894 28418
rect 10894 28366 10946 28418
rect 10946 28366 10948 28418
rect 10892 28364 10948 28366
rect 10556 28028 10612 28084
rect 11116 28028 11172 28084
rect 11228 29708 11284 29764
rect 10780 27858 10836 27860
rect 10780 27806 10782 27858
rect 10782 27806 10834 27858
rect 10834 27806 10836 27858
rect 10780 27804 10836 27806
rect 10556 27020 10612 27076
rect 10556 26514 10612 26516
rect 10556 26462 10558 26514
rect 10558 26462 10610 26514
rect 10610 26462 10612 26514
rect 10556 26460 10612 26462
rect 10556 26124 10612 26180
rect 11004 26402 11060 26404
rect 11004 26350 11006 26402
rect 11006 26350 11058 26402
rect 11058 26350 11060 26402
rect 11004 26348 11060 26350
rect 12460 32284 12516 32340
rect 12460 32060 12516 32116
rect 11900 30268 11956 30324
rect 12124 30828 12180 30884
rect 11788 30044 11844 30100
rect 11564 29932 11620 29988
rect 11900 29708 11956 29764
rect 12124 30098 12180 30100
rect 12124 30046 12126 30098
rect 12126 30046 12178 30098
rect 12178 30046 12180 30098
rect 12124 30044 12180 30046
rect 11788 29538 11844 29540
rect 11788 29486 11790 29538
rect 11790 29486 11842 29538
rect 11842 29486 11844 29538
rect 11788 29484 11844 29486
rect 11900 29372 11956 29428
rect 11340 28812 11396 28868
rect 12124 29372 12180 29428
rect 12460 29708 12516 29764
rect 12572 31106 12628 31108
rect 12572 31054 12574 31106
rect 12574 31054 12626 31106
rect 12626 31054 12628 31106
rect 12572 31052 12628 31054
rect 12908 33964 12964 34020
rect 13020 33404 13076 33460
rect 13356 36988 13412 37044
rect 13020 33122 13076 33124
rect 13020 33070 13022 33122
rect 13022 33070 13074 33122
rect 13074 33070 13076 33122
rect 13020 33068 13076 33070
rect 12796 32284 12852 32340
rect 13132 32562 13188 32564
rect 13132 32510 13134 32562
rect 13134 32510 13186 32562
rect 13186 32510 13188 32562
rect 13132 32508 13188 32510
rect 13132 31948 13188 32004
rect 13244 33628 13300 33684
rect 12908 31554 12964 31556
rect 12908 31502 12910 31554
rect 12910 31502 12962 31554
rect 12962 31502 12964 31554
rect 12908 31500 12964 31502
rect 13132 31276 13188 31332
rect 13692 37826 13748 37828
rect 13692 37774 13694 37826
rect 13694 37774 13746 37826
rect 13746 37774 13748 37826
rect 13692 37772 13748 37774
rect 13692 37212 13748 37268
rect 13580 36988 13636 37044
rect 14252 42140 14308 42196
rect 14028 41186 14084 41188
rect 14028 41134 14030 41186
rect 14030 41134 14082 41186
rect 14082 41134 14084 41186
rect 14028 41132 14084 41134
rect 14140 41020 14196 41076
rect 14364 40402 14420 40404
rect 14364 40350 14366 40402
rect 14366 40350 14418 40402
rect 14418 40350 14420 40402
rect 14364 40348 14420 40350
rect 14028 39004 14084 39060
rect 13916 38220 13972 38276
rect 14252 39228 14308 39284
rect 14140 38332 14196 38388
rect 13916 37826 13972 37828
rect 13916 37774 13918 37826
rect 13918 37774 13970 37826
rect 13970 37774 13972 37826
rect 13916 37772 13972 37774
rect 13916 37548 13972 37604
rect 14476 39452 14532 39508
rect 14476 38220 14532 38276
rect 14364 37548 14420 37604
rect 14028 36988 14084 37044
rect 13804 36428 13860 36484
rect 13692 36092 13748 36148
rect 14140 36706 14196 36708
rect 14140 36654 14142 36706
rect 14142 36654 14194 36706
rect 14194 36654 14196 36706
rect 14140 36652 14196 36654
rect 13468 35644 13524 35700
rect 13468 34914 13524 34916
rect 13468 34862 13470 34914
rect 13470 34862 13522 34914
rect 13522 34862 13524 34914
rect 13468 34860 13524 34862
rect 13580 34690 13636 34692
rect 13580 34638 13582 34690
rect 13582 34638 13634 34690
rect 13634 34638 13636 34690
rect 13580 34636 13636 34638
rect 13916 35868 13972 35924
rect 13916 34524 13972 34580
rect 14028 33628 14084 33684
rect 14140 35420 14196 35476
rect 14364 36482 14420 36484
rect 14364 36430 14366 36482
rect 14366 36430 14418 36482
rect 14418 36430 14420 36482
rect 14364 36428 14420 36430
rect 14476 34860 14532 34916
rect 14364 34636 14420 34692
rect 14252 34412 14308 34468
rect 14252 33516 14308 33572
rect 14812 44604 14868 44660
rect 15708 46396 15764 46452
rect 15820 46060 15876 46116
rect 15708 43932 15764 43988
rect 15260 43708 15316 43764
rect 15596 43708 15652 43764
rect 14924 41356 14980 41412
rect 15148 42588 15204 42644
rect 15036 41132 15092 41188
rect 14700 40012 14756 40068
rect 14700 39506 14756 39508
rect 14700 39454 14702 39506
rect 14702 39454 14754 39506
rect 14754 39454 14756 39506
rect 14700 39452 14756 39454
rect 15036 40012 15092 40068
rect 14812 39340 14868 39396
rect 15260 40460 15316 40516
rect 15036 39116 15092 39172
rect 15372 40012 15428 40068
rect 15708 40796 15764 40852
rect 15596 40348 15652 40404
rect 14812 38332 14868 38388
rect 15484 38834 15540 38836
rect 15484 38782 15486 38834
rect 15486 38782 15538 38834
rect 15538 38782 15540 38834
rect 15484 38780 15540 38782
rect 15036 37884 15092 37940
rect 15148 37324 15204 37380
rect 15708 39788 15764 39844
rect 15708 38332 15764 38388
rect 16044 48188 16100 48244
rect 16156 47404 16212 47460
rect 16044 47068 16100 47124
rect 17052 51548 17108 51604
rect 16828 51100 16884 51156
rect 16492 50428 16548 50484
rect 17724 51100 17780 51156
rect 17612 50428 17668 50484
rect 18060 52946 18116 52948
rect 18060 52894 18062 52946
rect 18062 52894 18114 52946
rect 18114 52894 18116 52946
rect 18060 52892 18116 52894
rect 18172 52834 18228 52836
rect 18172 52782 18174 52834
rect 18174 52782 18226 52834
rect 18226 52782 18228 52834
rect 18172 52780 18228 52782
rect 18396 54514 18452 54516
rect 18396 54462 18398 54514
rect 18398 54462 18450 54514
rect 18450 54462 18452 54514
rect 18396 54460 18452 54462
rect 18060 52220 18116 52276
rect 18396 52444 18452 52500
rect 18172 51996 18228 52052
rect 19068 52444 19124 52500
rect 20524 55410 20580 55412
rect 20524 55358 20526 55410
rect 20526 55358 20578 55410
rect 20578 55358 20580 55410
rect 20524 55356 20580 55358
rect 19836 54906 19892 54908
rect 19836 54854 19838 54906
rect 19838 54854 19890 54906
rect 19890 54854 19892 54906
rect 19836 54852 19892 54854
rect 19940 54906 19996 54908
rect 19940 54854 19942 54906
rect 19942 54854 19994 54906
rect 19994 54854 19996 54906
rect 19940 54852 19996 54854
rect 20044 54906 20100 54908
rect 20044 54854 20046 54906
rect 20046 54854 20098 54906
rect 20098 54854 20100 54906
rect 20044 54852 20100 54854
rect 19836 53338 19892 53340
rect 19836 53286 19838 53338
rect 19838 53286 19890 53338
rect 19890 53286 19892 53338
rect 19836 53284 19892 53286
rect 19940 53338 19996 53340
rect 19940 53286 19942 53338
rect 19942 53286 19994 53338
rect 19994 53286 19996 53338
rect 19940 53284 19996 53286
rect 20044 53338 20100 53340
rect 20044 53286 20046 53338
rect 20046 53286 20098 53338
rect 20098 53286 20100 53338
rect 20044 53284 20100 53286
rect 19180 52220 19236 52276
rect 19964 52780 20020 52836
rect 18620 52108 18676 52164
rect 20636 52162 20692 52164
rect 20636 52110 20638 52162
rect 20638 52110 20690 52162
rect 20690 52110 20692 52162
rect 20636 52108 20692 52110
rect 21084 52108 21140 52164
rect 19836 51770 19892 51772
rect 19836 51718 19838 51770
rect 19838 51718 19890 51770
rect 19890 51718 19892 51770
rect 19836 51716 19892 51718
rect 19940 51770 19996 51772
rect 19940 51718 19942 51770
rect 19942 51718 19994 51770
rect 19994 51718 19996 51770
rect 19940 51716 19996 51718
rect 20044 51770 20100 51772
rect 20044 51718 20046 51770
rect 20046 51718 20098 51770
rect 20098 51718 20100 51770
rect 20044 51716 20100 51718
rect 17948 50316 18004 50372
rect 17836 49868 17892 49924
rect 16492 48188 16548 48244
rect 18284 50370 18340 50372
rect 18284 50318 18286 50370
rect 18286 50318 18338 50370
rect 18338 50318 18340 50370
rect 18284 50316 18340 50318
rect 17612 48130 17668 48132
rect 17612 48078 17614 48130
rect 17614 48078 17666 48130
rect 17666 48078 17668 48130
rect 17612 48076 17668 48078
rect 18060 48076 18116 48132
rect 18396 49868 18452 49924
rect 19836 50202 19892 50204
rect 19836 50150 19838 50202
rect 19838 50150 19890 50202
rect 19890 50150 19892 50202
rect 19836 50148 19892 50150
rect 19940 50202 19996 50204
rect 19940 50150 19942 50202
rect 19942 50150 19994 50202
rect 19994 50150 19996 50202
rect 19940 50148 19996 50150
rect 20044 50202 20100 50204
rect 20044 50150 20046 50202
rect 20046 50150 20098 50202
rect 20098 50150 20100 50202
rect 20044 50148 20100 50150
rect 19068 48972 19124 49028
rect 20412 48914 20468 48916
rect 20412 48862 20414 48914
rect 20414 48862 20466 48914
rect 20466 48862 20468 48914
rect 20412 48860 20468 48862
rect 17164 47458 17220 47460
rect 17164 47406 17166 47458
rect 17166 47406 17218 47458
rect 17218 47406 17220 47458
rect 17164 47404 17220 47406
rect 18284 47852 18340 47908
rect 18620 48076 18676 48132
rect 18620 47740 18676 47796
rect 18508 47682 18564 47684
rect 18508 47630 18510 47682
rect 18510 47630 18562 47682
rect 18562 47630 18564 47682
rect 18508 47628 18564 47630
rect 18284 47458 18340 47460
rect 18284 47406 18286 47458
rect 18286 47406 18338 47458
rect 18338 47406 18340 47458
rect 18284 47404 18340 47406
rect 16380 46396 16436 46452
rect 16716 45890 16772 45892
rect 16716 45838 16718 45890
rect 16718 45838 16770 45890
rect 16770 45838 16772 45890
rect 16716 45836 16772 45838
rect 17388 45836 17444 45892
rect 16492 45724 16548 45780
rect 16268 44940 16324 44996
rect 17388 44828 17444 44884
rect 17500 44380 17556 44436
rect 16268 43932 16324 43988
rect 16156 40684 16212 40740
rect 15708 37996 15764 38052
rect 15708 37826 15764 37828
rect 15708 37774 15710 37826
rect 15710 37774 15762 37826
rect 15762 37774 15764 37826
rect 15708 37772 15764 37774
rect 14924 36652 14980 36708
rect 15036 35922 15092 35924
rect 15036 35870 15038 35922
rect 15038 35870 15090 35922
rect 15090 35870 15092 35922
rect 15036 35868 15092 35870
rect 14924 35308 14980 35364
rect 15372 35586 15428 35588
rect 15372 35534 15374 35586
rect 15374 35534 15426 35586
rect 15426 35534 15428 35586
rect 15372 35532 15428 35534
rect 15372 35308 15428 35364
rect 14700 34972 14756 35028
rect 14700 34636 14756 34692
rect 14812 34412 14868 34468
rect 14924 33964 14980 34020
rect 15036 34300 15092 34356
rect 14700 33852 14756 33908
rect 15596 34076 15652 34132
rect 14588 33516 14644 33572
rect 14028 33180 14084 33236
rect 13916 32674 13972 32676
rect 13916 32622 13918 32674
rect 13918 32622 13970 32674
rect 13970 32622 13972 32674
rect 13916 32620 13972 32622
rect 13580 32508 13636 32564
rect 13356 32060 13412 32116
rect 13356 31836 13412 31892
rect 13916 31724 13972 31780
rect 13468 31052 13524 31108
rect 13804 31276 13860 31332
rect 12236 28812 12292 28868
rect 11564 28082 11620 28084
rect 11564 28030 11566 28082
rect 11566 28030 11618 28082
rect 11618 28030 11620 28082
rect 11564 28028 11620 28030
rect 12236 28028 12292 28084
rect 12124 27858 12180 27860
rect 12124 27806 12126 27858
rect 12126 27806 12178 27858
rect 12178 27806 12180 27858
rect 12124 27804 12180 27806
rect 12348 27244 12404 27300
rect 12236 27074 12292 27076
rect 12236 27022 12238 27074
rect 12238 27022 12290 27074
rect 12290 27022 12292 27074
rect 12236 27020 12292 27022
rect 11788 26796 11844 26852
rect 11452 26572 11508 26628
rect 11004 25900 11060 25956
rect 11004 25506 11060 25508
rect 11004 25454 11006 25506
rect 11006 25454 11058 25506
rect 11058 25454 11060 25506
rect 11004 25452 11060 25454
rect 10444 25340 10500 25396
rect 10780 25394 10836 25396
rect 10780 25342 10782 25394
rect 10782 25342 10834 25394
rect 10834 25342 10836 25394
rect 10780 25340 10836 25342
rect 12012 26572 12068 26628
rect 11900 26290 11956 26292
rect 11900 26238 11902 26290
rect 11902 26238 11954 26290
rect 11954 26238 11956 26290
rect 11900 26236 11956 26238
rect 11900 25506 11956 25508
rect 11900 25454 11902 25506
rect 11902 25454 11954 25506
rect 11954 25454 11956 25506
rect 11900 25452 11956 25454
rect 11676 24946 11732 24948
rect 11676 24894 11678 24946
rect 11678 24894 11730 24946
rect 11730 24894 11732 24946
rect 11676 24892 11732 24894
rect 12684 29986 12740 29988
rect 12684 29934 12686 29986
rect 12686 29934 12738 29986
rect 12738 29934 12740 29986
rect 12684 29932 12740 29934
rect 12684 29260 12740 29316
rect 12684 28754 12740 28756
rect 12684 28702 12686 28754
rect 12686 28702 12738 28754
rect 12738 28702 12740 28754
rect 12684 28700 12740 28702
rect 12572 28476 12628 28532
rect 12684 27804 12740 27860
rect 13020 30716 13076 30772
rect 13692 30044 13748 30100
rect 13580 29820 13636 29876
rect 13356 29708 13412 29764
rect 13356 28700 13412 28756
rect 14028 31948 14084 32004
rect 14252 32674 14308 32676
rect 14252 32622 14254 32674
rect 14254 32622 14306 32674
rect 14306 32622 14308 32674
rect 14252 32620 14308 32622
rect 14588 32620 14644 32676
rect 15036 33122 15092 33124
rect 15036 33070 15038 33122
rect 15038 33070 15090 33122
rect 15090 33070 15092 33122
rect 15036 33068 15092 33070
rect 14252 31052 14308 31108
rect 14476 31052 14532 31108
rect 14140 30940 14196 30996
rect 14140 30604 14196 30660
rect 14812 31778 14868 31780
rect 14812 31726 14814 31778
rect 14814 31726 14866 31778
rect 14866 31726 14868 31778
rect 14812 31724 14868 31726
rect 14588 30380 14644 30436
rect 13692 29260 13748 29316
rect 15036 32844 15092 32900
rect 15260 31948 15316 32004
rect 15260 31612 15316 31668
rect 15484 33458 15540 33460
rect 15484 33406 15486 33458
rect 15486 33406 15538 33458
rect 15538 33406 15540 33458
rect 15484 33404 15540 33406
rect 15372 31164 15428 31220
rect 15484 31106 15540 31108
rect 15484 31054 15486 31106
rect 15486 31054 15538 31106
rect 15538 31054 15540 31106
rect 15484 31052 15540 31054
rect 15036 30604 15092 30660
rect 15260 30940 15316 30996
rect 14924 30044 14980 30100
rect 15148 29932 15204 29988
rect 14812 29372 14868 29428
rect 16604 44322 16660 44324
rect 16604 44270 16606 44322
rect 16606 44270 16658 44322
rect 16658 44270 16660 44322
rect 16604 44268 16660 44270
rect 16828 44322 16884 44324
rect 16828 44270 16830 44322
rect 16830 44270 16882 44322
rect 16882 44270 16884 44322
rect 16828 44268 16884 44270
rect 16380 43708 16436 43764
rect 16604 43484 16660 43540
rect 16380 41132 16436 41188
rect 16380 39788 16436 39844
rect 16716 42700 16772 42756
rect 17388 44210 17444 44212
rect 17388 44158 17390 44210
rect 17390 44158 17442 44210
rect 17442 44158 17444 44210
rect 17388 44156 17444 44158
rect 17276 44098 17332 44100
rect 17276 44046 17278 44098
rect 17278 44046 17330 44098
rect 17330 44046 17332 44098
rect 17276 44044 17332 44046
rect 18172 47068 18228 47124
rect 17836 45778 17892 45780
rect 17836 45726 17838 45778
rect 17838 45726 17890 45778
rect 17890 45726 17892 45778
rect 17836 45724 17892 45726
rect 17724 45052 17780 45108
rect 17724 44044 17780 44100
rect 17500 43762 17556 43764
rect 17500 43710 17502 43762
rect 17502 43710 17554 43762
rect 17554 43710 17556 43762
rect 17500 43708 17556 43710
rect 17612 43650 17668 43652
rect 17612 43598 17614 43650
rect 17614 43598 17666 43650
rect 17666 43598 17668 43650
rect 17612 43596 17668 43598
rect 17052 42700 17108 42756
rect 17612 42754 17668 42756
rect 17612 42702 17614 42754
rect 17614 42702 17666 42754
rect 17666 42702 17668 42754
rect 17612 42700 17668 42702
rect 16604 41970 16660 41972
rect 16604 41918 16606 41970
rect 16606 41918 16658 41970
rect 16658 41918 16660 41970
rect 16604 41916 16660 41918
rect 16604 40012 16660 40068
rect 18060 42476 18116 42532
rect 17836 42364 17892 42420
rect 18060 42028 18116 42084
rect 17948 41916 18004 41972
rect 16380 38220 16436 38276
rect 16492 38332 16548 38388
rect 16268 37996 16324 38052
rect 16380 37826 16436 37828
rect 16380 37774 16382 37826
rect 16382 37774 16434 37826
rect 16434 37774 16436 37826
rect 16380 37772 16436 37774
rect 16156 37324 16212 37380
rect 16268 37266 16324 37268
rect 16268 37214 16270 37266
rect 16270 37214 16322 37266
rect 16322 37214 16324 37266
rect 16268 37212 16324 37214
rect 16492 37548 16548 37604
rect 16492 37378 16548 37380
rect 16492 37326 16494 37378
rect 16494 37326 16546 37378
rect 16546 37326 16548 37378
rect 16492 37324 16548 37326
rect 16380 36204 16436 36260
rect 16044 35868 16100 35924
rect 16268 35532 16324 35588
rect 15932 34972 15988 35028
rect 15932 33180 15988 33236
rect 16156 33180 16212 33236
rect 16940 38780 16996 38836
rect 17612 41186 17668 41188
rect 17612 41134 17614 41186
rect 17614 41134 17666 41186
rect 17666 41134 17668 41186
rect 17612 41132 17668 41134
rect 17500 40684 17556 40740
rect 17500 40460 17556 40516
rect 17724 40124 17780 40180
rect 17388 39676 17444 39732
rect 17276 37436 17332 37492
rect 17836 38050 17892 38052
rect 17836 37998 17838 38050
rect 17838 37998 17890 38050
rect 17890 37998 17892 38050
rect 17836 37996 17892 37998
rect 17724 37938 17780 37940
rect 17724 37886 17726 37938
rect 17726 37886 17778 37938
rect 17778 37886 17780 37938
rect 17724 37884 17780 37886
rect 17388 37212 17444 37268
rect 16940 34914 16996 34916
rect 16940 34862 16942 34914
rect 16942 34862 16994 34914
rect 16994 34862 16996 34914
rect 16940 34860 16996 34862
rect 16828 34802 16884 34804
rect 16828 34750 16830 34802
rect 16830 34750 16882 34802
rect 16882 34750 16884 34802
rect 16828 34748 16884 34750
rect 17052 34188 17108 34244
rect 16716 34130 16772 34132
rect 16716 34078 16718 34130
rect 16718 34078 16770 34130
rect 16770 34078 16772 34130
rect 16716 34076 16772 34078
rect 16604 33628 16660 33684
rect 16940 33740 16996 33796
rect 17052 33628 17108 33684
rect 17500 37548 17556 37604
rect 17500 36370 17556 36372
rect 17500 36318 17502 36370
rect 17502 36318 17554 36370
rect 17554 36318 17556 36370
rect 17500 36316 17556 36318
rect 18172 41970 18228 41972
rect 18172 41918 18174 41970
rect 18174 41918 18226 41970
rect 18226 41918 18228 41970
rect 18172 41916 18228 41918
rect 18620 47068 18676 47124
rect 18620 44492 18676 44548
rect 19180 48076 19236 48132
rect 18956 47852 19012 47908
rect 18956 47628 19012 47684
rect 18732 44156 18788 44212
rect 19836 48634 19892 48636
rect 19836 48582 19838 48634
rect 19838 48582 19890 48634
rect 19890 48582 19892 48634
rect 19836 48580 19892 48582
rect 19940 48634 19996 48636
rect 19940 48582 19942 48634
rect 19942 48582 19994 48634
rect 19994 48582 19996 48634
rect 19940 48580 19996 48582
rect 20044 48634 20100 48636
rect 20044 48582 20046 48634
rect 20046 48582 20098 48634
rect 20098 48582 20100 48634
rect 20044 48580 20100 48582
rect 19628 48354 19684 48356
rect 19628 48302 19630 48354
rect 19630 48302 19682 48354
rect 19682 48302 19684 48354
rect 19628 48300 19684 48302
rect 20524 48188 20580 48244
rect 20076 47628 20132 47684
rect 20076 47458 20132 47460
rect 20076 47406 20078 47458
rect 20078 47406 20130 47458
rect 20130 47406 20132 47458
rect 20076 47404 20132 47406
rect 19836 47066 19892 47068
rect 19836 47014 19838 47066
rect 19838 47014 19890 47066
rect 19890 47014 19892 47066
rect 19836 47012 19892 47014
rect 19940 47066 19996 47068
rect 19940 47014 19942 47066
rect 19942 47014 19994 47066
rect 19994 47014 19996 47066
rect 19940 47012 19996 47014
rect 20044 47066 20100 47068
rect 20044 47014 20046 47066
rect 20046 47014 20098 47066
rect 20098 47014 20100 47066
rect 20044 47012 20100 47014
rect 19628 46508 19684 46564
rect 20076 46620 20132 46676
rect 18620 43538 18676 43540
rect 18620 43486 18622 43538
rect 18622 43486 18674 43538
rect 18674 43486 18676 43538
rect 18620 43484 18676 43486
rect 20300 45836 20356 45892
rect 19628 45500 19684 45556
rect 19836 45498 19892 45500
rect 19836 45446 19838 45498
rect 19838 45446 19890 45498
rect 19890 45446 19892 45498
rect 19836 45444 19892 45446
rect 19940 45498 19996 45500
rect 19940 45446 19942 45498
rect 19942 45446 19994 45498
rect 19994 45446 19996 45498
rect 19940 45444 19996 45446
rect 20044 45498 20100 45500
rect 20044 45446 20046 45498
rect 20046 45446 20098 45498
rect 20098 45446 20100 45498
rect 20044 45444 20100 45446
rect 20188 45500 20244 45556
rect 20300 44994 20356 44996
rect 20300 44942 20302 44994
rect 20302 44942 20354 44994
rect 20354 44942 20356 44994
rect 20300 44940 20356 44942
rect 19964 44604 20020 44660
rect 19628 44380 19684 44436
rect 19852 44210 19908 44212
rect 19852 44158 19854 44210
rect 19854 44158 19906 44210
rect 19906 44158 19908 44210
rect 19852 44156 19908 44158
rect 19068 43596 19124 43652
rect 19292 44044 19348 44100
rect 18732 42924 18788 42980
rect 18732 42588 18788 42644
rect 18284 40684 18340 40740
rect 18172 40626 18228 40628
rect 18172 40574 18174 40626
rect 18174 40574 18226 40626
rect 18226 40574 18228 40626
rect 18172 40572 18228 40574
rect 18508 40290 18564 40292
rect 18508 40238 18510 40290
rect 18510 40238 18562 40290
rect 18562 40238 18564 40290
rect 18508 40236 18564 40238
rect 18172 39506 18228 39508
rect 18172 39454 18174 39506
rect 18174 39454 18226 39506
rect 18226 39454 18228 39506
rect 18172 39452 18228 39454
rect 18844 41746 18900 41748
rect 18844 41694 18846 41746
rect 18846 41694 18898 41746
rect 18898 41694 18900 41746
rect 18844 41692 18900 41694
rect 18732 40572 18788 40628
rect 18172 38892 18228 38948
rect 18284 37548 18340 37604
rect 18956 39228 19012 39284
rect 18508 38050 18564 38052
rect 18508 37998 18510 38050
rect 18510 37998 18562 38050
rect 18562 37998 18564 38050
rect 18508 37996 18564 37998
rect 18396 37436 18452 37492
rect 18284 37378 18340 37380
rect 18284 37326 18286 37378
rect 18286 37326 18338 37378
rect 18338 37326 18340 37378
rect 18284 37324 18340 37326
rect 17836 37212 17892 37268
rect 18396 36764 18452 36820
rect 18060 36652 18116 36708
rect 18956 37772 19012 37828
rect 19068 37884 19124 37940
rect 19180 37660 19236 37716
rect 19180 37490 19236 37492
rect 19180 37438 19182 37490
rect 19182 37438 19234 37490
rect 19234 37438 19236 37490
rect 19180 37436 19236 37438
rect 18508 36652 18564 36708
rect 18620 37100 18676 37156
rect 17948 36428 18004 36484
rect 17836 36258 17892 36260
rect 17836 36206 17838 36258
rect 17838 36206 17890 36258
rect 17890 36206 17892 36258
rect 17836 36204 17892 36206
rect 18172 36092 18228 36148
rect 17724 35810 17780 35812
rect 17724 35758 17726 35810
rect 17726 35758 17778 35810
rect 17778 35758 17780 35810
rect 17724 35756 17780 35758
rect 17948 34412 18004 34468
rect 17612 34300 17668 34356
rect 17500 34242 17556 34244
rect 17500 34190 17502 34242
rect 17502 34190 17554 34242
rect 17554 34190 17556 34242
rect 17500 34188 17556 34190
rect 17612 33964 17668 34020
rect 17388 33516 17444 33572
rect 16940 33068 16996 33124
rect 17164 33068 17220 33124
rect 16156 31948 16212 32004
rect 15708 31052 15764 31108
rect 14364 28700 14420 28756
rect 13244 28476 13300 28532
rect 13244 27804 13300 27860
rect 13580 27074 13636 27076
rect 13580 27022 13582 27074
rect 13582 27022 13634 27074
rect 13634 27022 13636 27074
rect 13580 27020 13636 27022
rect 12572 25394 12628 25396
rect 12572 25342 12574 25394
rect 12574 25342 12626 25394
rect 12626 25342 12628 25394
rect 12572 25340 12628 25342
rect 12460 25228 12516 25284
rect 12348 24892 12404 24948
rect 11340 24108 11396 24164
rect 11676 24668 11732 24724
rect 10332 23324 10388 23380
rect 13692 26572 13748 26628
rect 12796 26514 12852 26516
rect 12796 26462 12798 26514
rect 12798 26462 12850 26514
rect 12850 26462 12852 26514
rect 12796 26460 12852 26462
rect 13244 26514 13300 26516
rect 13244 26462 13246 26514
rect 13246 26462 13298 26514
rect 13298 26462 13300 26514
rect 13244 26460 13300 26462
rect 15260 28700 15316 28756
rect 14700 28530 14756 28532
rect 14700 28478 14702 28530
rect 14702 28478 14754 28530
rect 14754 28478 14756 28530
rect 14700 28476 14756 28478
rect 14140 28028 14196 28084
rect 14252 27692 14308 27748
rect 13916 26348 13972 26404
rect 13580 26236 13636 26292
rect 12908 24220 12964 24276
rect 13468 25282 13524 25284
rect 13468 25230 13470 25282
rect 13470 25230 13522 25282
rect 13522 25230 13524 25282
rect 13468 25228 13524 25230
rect 13356 24780 13412 24836
rect 14140 25788 14196 25844
rect 13916 25228 13972 25284
rect 14028 25116 14084 25172
rect 14476 27244 14532 27300
rect 14924 28530 14980 28532
rect 14924 28478 14926 28530
rect 14926 28478 14978 28530
rect 14978 28478 14980 28530
rect 14924 28476 14980 28478
rect 15148 27916 15204 27972
rect 15372 28364 15428 28420
rect 14812 27132 14868 27188
rect 16156 31164 16212 31220
rect 16044 30940 16100 30996
rect 16044 30492 16100 30548
rect 16268 30940 16324 30996
rect 16492 32450 16548 32452
rect 16492 32398 16494 32450
rect 16494 32398 16546 32450
rect 16546 32398 16548 32450
rect 16492 32396 16548 32398
rect 16828 32562 16884 32564
rect 16828 32510 16830 32562
rect 16830 32510 16882 32562
rect 16882 32510 16884 32562
rect 16828 32508 16884 32510
rect 16604 32284 16660 32340
rect 16156 30156 16212 30212
rect 16828 32284 16884 32340
rect 15596 28028 15652 28084
rect 15484 27858 15540 27860
rect 15484 27806 15486 27858
rect 15486 27806 15538 27858
rect 15538 27806 15540 27858
rect 15484 27804 15540 27806
rect 15148 26962 15204 26964
rect 15148 26910 15150 26962
rect 15150 26910 15202 26962
rect 15202 26910 15204 26962
rect 15148 26908 15204 26910
rect 15820 27580 15876 27636
rect 16044 28364 16100 28420
rect 15708 27132 15764 27188
rect 16716 31948 16772 32004
rect 17052 32002 17108 32004
rect 17052 31950 17054 32002
rect 17054 31950 17106 32002
rect 17106 31950 17108 32002
rect 17052 31948 17108 31950
rect 16604 31778 16660 31780
rect 16604 31726 16606 31778
rect 16606 31726 16658 31778
rect 16658 31726 16660 31778
rect 16604 31724 16660 31726
rect 16492 30044 16548 30100
rect 17052 31276 17108 31332
rect 17276 31276 17332 31332
rect 16828 30994 16884 30996
rect 16828 30942 16830 30994
rect 16830 30942 16882 30994
rect 16882 30942 16884 30994
rect 16828 30940 16884 30942
rect 17164 30828 17220 30884
rect 17500 33346 17556 33348
rect 17500 33294 17502 33346
rect 17502 33294 17554 33346
rect 17554 33294 17556 33346
rect 17500 33292 17556 33294
rect 17724 33852 17780 33908
rect 17276 30044 17332 30100
rect 15036 26796 15092 26852
rect 15708 26796 15764 26852
rect 15596 26684 15652 26740
rect 15036 26514 15092 26516
rect 15036 26462 15038 26514
rect 15038 26462 15090 26514
rect 15090 26462 15092 26514
rect 15036 26460 15092 26462
rect 15260 26572 15316 26628
rect 14476 25788 14532 25844
rect 14700 25452 14756 25508
rect 15372 26460 15428 26516
rect 15708 26236 15764 26292
rect 15596 25340 15652 25396
rect 14252 24780 14308 24836
rect 16268 27468 16324 27524
rect 16156 26348 16212 26404
rect 16268 27244 16324 27300
rect 16044 26290 16100 26292
rect 16044 26238 16046 26290
rect 16046 26238 16098 26290
rect 16098 26238 16100 26290
rect 16044 26236 16100 26238
rect 16716 28754 16772 28756
rect 16716 28702 16718 28754
rect 16718 28702 16770 28754
rect 16770 28702 16772 28754
rect 16716 28700 16772 28702
rect 16716 28476 16772 28532
rect 16716 27970 16772 27972
rect 16716 27918 16718 27970
rect 16718 27918 16770 27970
rect 16770 27918 16772 27970
rect 16716 27916 16772 27918
rect 16380 26796 16436 26852
rect 16716 27634 16772 27636
rect 16716 27582 16718 27634
rect 16718 27582 16770 27634
rect 16770 27582 16772 27634
rect 16716 27580 16772 27582
rect 17164 27244 17220 27300
rect 16604 26850 16660 26852
rect 16604 26798 16606 26850
rect 16606 26798 16658 26850
rect 16658 26798 16660 26850
rect 16604 26796 16660 26798
rect 16940 26796 16996 26852
rect 15932 25900 15988 25956
rect 16380 26124 16436 26180
rect 15820 25676 15876 25732
rect 16268 25676 16324 25732
rect 16044 25506 16100 25508
rect 16044 25454 16046 25506
rect 16046 25454 16098 25506
rect 16098 25454 16100 25506
rect 16044 25452 16100 25454
rect 16156 25340 16212 25396
rect 14700 24220 14756 24276
rect 15708 24108 15764 24164
rect 15148 24050 15204 24052
rect 15148 23998 15150 24050
rect 15150 23998 15202 24050
rect 15202 23998 15204 24050
rect 15148 23996 15204 23998
rect 15484 23938 15540 23940
rect 15484 23886 15486 23938
rect 15486 23886 15538 23938
rect 15538 23886 15540 23938
rect 15484 23884 15540 23886
rect 15820 23772 15876 23828
rect 15820 23266 15876 23268
rect 15820 23214 15822 23266
rect 15822 23214 15874 23266
rect 15874 23214 15876 23266
rect 15820 23212 15876 23214
rect 15148 22652 15204 22708
rect 16492 24722 16548 24724
rect 16492 24670 16494 24722
rect 16494 24670 16546 24722
rect 16546 24670 16548 24722
rect 16492 24668 16548 24670
rect 16716 25564 16772 25620
rect 16940 26124 16996 26180
rect 16828 25452 16884 25508
rect 16716 24668 16772 24724
rect 17724 32562 17780 32564
rect 17724 32510 17726 32562
rect 17726 32510 17778 32562
rect 17778 32510 17780 32562
rect 17724 32508 17780 32510
rect 17948 33740 18004 33796
rect 18060 33964 18116 34020
rect 17948 32956 18004 33012
rect 17948 32508 18004 32564
rect 18060 32450 18116 32452
rect 18060 32398 18062 32450
rect 18062 32398 18114 32450
rect 18114 32398 18116 32450
rect 18060 32396 18116 32398
rect 18284 34748 18340 34804
rect 18396 36204 18452 36260
rect 18620 36204 18676 36260
rect 19836 43930 19892 43932
rect 19836 43878 19838 43930
rect 19838 43878 19890 43930
rect 19890 43878 19892 43930
rect 19836 43876 19892 43878
rect 19940 43930 19996 43932
rect 19940 43878 19942 43930
rect 19942 43878 19994 43930
rect 19994 43878 19996 43930
rect 19940 43876 19996 43878
rect 20044 43930 20100 43932
rect 20044 43878 20046 43930
rect 20046 43878 20098 43930
rect 20098 43878 20100 43930
rect 20044 43876 20100 43878
rect 19836 42362 19892 42364
rect 19836 42310 19838 42362
rect 19838 42310 19890 42362
rect 19890 42310 19892 42362
rect 19836 42308 19892 42310
rect 19940 42362 19996 42364
rect 19940 42310 19942 42362
rect 19942 42310 19994 42362
rect 19994 42310 19996 42362
rect 19940 42308 19996 42310
rect 20044 42362 20100 42364
rect 20044 42310 20046 42362
rect 20046 42310 20098 42362
rect 20098 42310 20100 42362
rect 20044 42308 20100 42310
rect 20188 41970 20244 41972
rect 20188 41918 20190 41970
rect 20190 41918 20242 41970
rect 20242 41918 20244 41970
rect 20188 41916 20244 41918
rect 19516 41692 19572 41748
rect 19516 41132 19572 41188
rect 19852 41580 19908 41636
rect 20188 41356 20244 41412
rect 19852 41074 19908 41076
rect 19852 41022 19854 41074
rect 19854 41022 19906 41074
rect 19906 41022 19908 41074
rect 19852 41020 19908 41022
rect 19836 40794 19892 40796
rect 19836 40742 19838 40794
rect 19838 40742 19890 40794
rect 19890 40742 19892 40794
rect 19836 40740 19892 40742
rect 19940 40794 19996 40796
rect 19940 40742 19942 40794
rect 19942 40742 19994 40794
rect 19994 40742 19996 40794
rect 19940 40740 19996 40742
rect 20044 40794 20100 40796
rect 20044 40742 20046 40794
rect 20046 40742 20098 40794
rect 20098 40742 20100 40794
rect 20044 40740 20100 40742
rect 21420 55298 21476 55300
rect 21420 55246 21422 55298
rect 21422 55246 21474 55298
rect 21474 55246 21476 55298
rect 21420 55244 21476 55246
rect 23212 55356 23268 55412
rect 22876 54460 22932 54516
rect 21756 53676 21812 53732
rect 22428 53730 22484 53732
rect 22428 53678 22430 53730
rect 22430 53678 22482 53730
rect 22482 53678 22484 53730
rect 22428 53676 22484 53678
rect 22652 53730 22708 53732
rect 22652 53678 22654 53730
rect 22654 53678 22706 53730
rect 22706 53678 22708 53730
rect 22652 53676 22708 53678
rect 22316 53618 22372 53620
rect 22316 53566 22318 53618
rect 22318 53566 22370 53618
rect 22370 53566 22372 53618
rect 22316 53564 22372 53566
rect 21980 53506 22036 53508
rect 21980 53454 21982 53506
rect 21982 53454 22034 53506
rect 22034 53454 22036 53506
rect 21980 53452 22036 53454
rect 22652 53452 22708 53508
rect 22876 53788 22932 53844
rect 22764 53058 22820 53060
rect 22764 53006 22766 53058
rect 22766 53006 22818 53058
rect 22818 53006 22820 53058
rect 22764 53004 22820 53006
rect 21756 52780 21812 52836
rect 22540 52834 22596 52836
rect 22540 52782 22542 52834
rect 22542 52782 22594 52834
rect 22594 52782 22596 52834
rect 22540 52780 22596 52782
rect 22428 50764 22484 50820
rect 21868 50594 21924 50596
rect 21868 50542 21870 50594
rect 21870 50542 21922 50594
rect 21922 50542 21924 50594
rect 21868 50540 21924 50542
rect 22988 50652 23044 50708
rect 23100 52220 23156 52276
rect 22204 49868 22260 49924
rect 21868 49026 21924 49028
rect 21868 48974 21870 49026
rect 21870 48974 21922 49026
rect 21922 48974 21924 49026
rect 21868 48972 21924 48974
rect 21644 48242 21700 48244
rect 21644 48190 21646 48242
rect 21646 48190 21698 48242
rect 21698 48190 21700 48242
rect 21644 48188 21700 48190
rect 27916 56028 27972 56084
rect 28588 56082 28644 56084
rect 28588 56030 28590 56082
rect 28590 56030 28642 56082
rect 28642 56030 28644 56082
rect 28588 56028 28644 56030
rect 30492 55804 30548 55860
rect 29260 55298 29316 55300
rect 29260 55246 29262 55298
rect 29262 55246 29314 55298
rect 29314 55246 29316 55298
rect 29260 55244 29316 55246
rect 23436 54460 23492 54516
rect 23660 53842 23716 53844
rect 23660 53790 23662 53842
rect 23662 53790 23714 53842
rect 23714 53790 23716 53842
rect 23660 53788 23716 53790
rect 24892 54348 24948 54404
rect 23548 52892 23604 52948
rect 23996 53004 24052 53060
rect 23660 50706 23716 50708
rect 23660 50654 23662 50706
rect 23662 50654 23714 50706
rect 23714 50654 23716 50706
rect 23660 50652 23716 50654
rect 23548 50482 23604 50484
rect 23548 50430 23550 50482
rect 23550 50430 23602 50482
rect 23602 50430 23604 50482
rect 23548 50428 23604 50430
rect 24108 50540 24164 50596
rect 23772 49868 23828 49924
rect 24556 53564 24612 53620
rect 25228 53618 25284 53620
rect 25228 53566 25230 53618
rect 25230 53566 25282 53618
rect 25282 53566 25284 53618
rect 25228 53564 25284 53566
rect 25004 53452 25060 53508
rect 24892 52556 24948 52612
rect 25228 52108 25284 52164
rect 26012 54402 26068 54404
rect 26012 54350 26014 54402
rect 26014 54350 26066 54402
rect 26066 54350 26068 54402
rect 26012 54348 26068 54350
rect 29148 54684 29204 54740
rect 28812 54514 28868 54516
rect 28812 54462 28814 54514
rect 28814 54462 28866 54514
rect 28866 54462 28868 54514
rect 28812 54460 28868 54462
rect 27580 54348 27636 54404
rect 26572 53788 26628 53844
rect 26348 53618 26404 53620
rect 26348 53566 26350 53618
rect 26350 53566 26402 53618
rect 26402 53566 26404 53618
rect 26348 53564 26404 53566
rect 25676 53506 25732 53508
rect 25676 53454 25678 53506
rect 25678 53454 25730 53506
rect 25730 53454 25732 53506
rect 25676 53452 25732 53454
rect 25452 53004 25508 53060
rect 25452 52444 25508 52500
rect 25452 51996 25508 52052
rect 28140 53788 28196 53844
rect 29148 54236 29204 54292
rect 30044 54514 30100 54516
rect 30044 54462 30046 54514
rect 30046 54462 30098 54514
rect 30098 54462 30100 54514
rect 30044 54460 30100 54462
rect 27580 53676 27636 53732
rect 26124 52946 26180 52948
rect 26124 52894 26126 52946
rect 26126 52894 26178 52946
rect 26178 52894 26180 52946
rect 26124 52892 26180 52894
rect 25900 51212 25956 51268
rect 24444 50594 24500 50596
rect 24444 50542 24446 50594
rect 24446 50542 24498 50594
rect 24498 50542 24500 50594
rect 24444 50540 24500 50542
rect 26012 50540 26068 50596
rect 26236 50764 26292 50820
rect 24556 50428 24612 50484
rect 29260 53452 29316 53508
rect 26684 53058 26740 53060
rect 26684 53006 26686 53058
rect 26686 53006 26738 53058
rect 26738 53006 26740 53058
rect 26684 53004 26740 53006
rect 31836 54626 31892 54628
rect 31836 54574 31838 54626
rect 31838 54574 31890 54626
rect 31890 54574 31892 54626
rect 31836 54572 31892 54574
rect 30380 53788 30436 53844
rect 30268 53452 30324 53508
rect 30044 53058 30100 53060
rect 30044 53006 30046 53058
rect 30046 53006 30098 53058
rect 30098 53006 30100 53058
rect 30044 53004 30100 53006
rect 27020 52780 27076 52836
rect 27468 52834 27524 52836
rect 27468 52782 27470 52834
rect 27470 52782 27522 52834
rect 27522 52782 27524 52834
rect 27468 52780 27524 52782
rect 28476 52780 28532 52836
rect 27244 52220 27300 52276
rect 26796 51996 26852 52052
rect 26796 50764 26852 50820
rect 26908 51324 26964 51380
rect 26796 50594 26852 50596
rect 26796 50542 26798 50594
rect 26798 50542 26850 50594
rect 26850 50542 26852 50594
rect 26796 50540 26852 50542
rect 22428 48300 22484 48356
rect 22204 48188 22260 48244
rect 22428 47964 22484 48020
rect 21980 47852 22036 47908
rect 22540 47852 22596 47908
rect 22876 48636 22932 48692
rect 23212 48412 23268 48468
rect 23884 48412 23940 48468
rect 22876 48188 22932 48244
rect 21308 46620 21364 46676
rect 21084 45724 21140 45780
rect 20524 44380 20580 44436
rect 20748 45276 20804 45332
rect 20860 44940 20916 44996
rect 20972 44492 21028 44548
rect 20748 44322 20804 44324
rect 20748 44270 20750 44322
rect 20750 44270 20802 44322
rect 20802 44270 20804 44322
rect 20748 44268 20804 44270
rect 20748 42364 20804 42420
rect 21196 45388 21252 45444
rect 20636 41580 20692 41636
rect 20524 41074 20580 41076
rect 20524 41022 20526 41074
rect 20526 41022 20578 41074
rect 20578 41022 20580 41074
rect 20524 41020 20580 41022
rect 20188 40572 20244 40628
rect 19516 39900 19572 39956
rect 19404 39340 19460 39396
rect 20076 39788 20132 39844
rect 20188 39340 20244 39396
rect 19836 39226 19892 39228
rect 19836 39174 19838 39226
rect 19838 39174 19890 39226
rect 19890 39174 19892 39226
rect 19836 39172 19892 39174
rect 19940 39226 19996 39228
rect 19940 39174 19942 39226
rect 19942 39174 19994 39226
rect 19994 39174 19996 39226
rect 19940 39172 19996 39174
rect 20044 39226 20100 39228
rect 20044 39174 20046 39226
rect 20046 39174 20098 39226
rect 20098 39174 20100 39226
rect 20044 39172 20100 39174
rect 19740 38220 19796 38276
rect 19964 38050 20020 38052
rect 19964 37998 19966 38050
rect 19966 37998 20018 38050
rect 20018 37998 20020 38050
rect 19964 37996 20020 37998
rect 19740 37938 19796 37940
rect 19740 37886 19742 37938
rect 19742 37886 19794 37938
rect 19794 37886 19796 37938
rect 19740 37884 19796 37886
rect 19628 37772 19684 37828
rect 19404 37490 19460 37492
rect 19404 37438 19406 37490
rect 19406 37438 19458 37490
rect 19458 37438 19460 37490
rect 19404 37436 19460 37438
rect 19404 36876 19460 36932
rect 18956 36258 19012 36260
rect 18956 36206 18958 36258
rect 18958 36206 19010 36258
rect 19010 36206 19012 36258
rect 18956 36204 19012 36206
rect 18844 35756 18900 35812
rect 18620 35420 18676 35476
rect 18508 35084 18564 35140
rect 18844 35196 18900 35252
rect 18508 34860 18564 34916
rect 18844 34802 18900 34804
rect 18844 34750 18846 34802
rect 18846 34750 18898 34802
rect 18898 34750 18900 34802
rect 18844 34748 18900 34750
rect 19180 36540 19236 36596
rect 19180 36092 19236 36148
rect 19292 35810 19348 35812
rect 19292 35758 19294 35810
rect 19294 35758 19346 35810
rect 19346 35758 19348 35810
rect 19292 35756 19348 35758
rect 19180 35196 19236 35252
rect 19068 34690 19124 34692
rect 19068 34638 19070 34690
rect 19070 34638 19122 34690
rect 19122 34638 19124 34690
rect 19068 34636 19124 34638
rect 18396 33852 18452 33908
rect 18284 33404 18340 33460
rect 18284 33234 18340 33236
rect 18284 33182 18286 33234
rect 18286 33182 18338 33234
rect 18338 33182 18340 33234
rect 18284 33180 18340 33182
rect 18284 32956 18340 33012
rect 19068 34130 19124 34132
rect 19068 34078 19070 34130
rect 19070 34078 19122 34130
rect 19122 34078 19124 34130
rect 19068 34076 19124 34078
rect 19836 37658 19892 37660
rect 19836 37606 19838 37658
rect 19838 37606 19890 37658
rect 19890 37606 19892 37658
rect 19836 37604 19892 37606
rect 19940 37658 19996 37660
rect 19940 37606 19942 37658
rect 19942 37606 19994 37658
rect 19994 37606 19996 37658
rect 19940 37604 19996 37606
rect 20044 37658 20100 37660
rect 20044 37606 20046 37658
rect 20046 37606 20098 37658
rect 20098 37606 20100 37658
rect 20044 37604 20100 37606
rect 21756 46508 21812 46564
rect 21420 45836 21476 45892
rect 21420 45500 21476 45556
rect 21644 44604 21700 44660
rect 21756 44492 21812 44548
rect 22540 46844 22596 46900
rect 21868 44156 21924 44212
rect 21084 42812 21140 42868
rect 21756 43260 21812 43316
rect 20972 41970 21028 41972
rect 20972 41918 20974 41970
rect 20974 41918 21026 41970
rect 21026 41918 21028 41970
rect 20972 41916 21028 41918
rect 20860 41580 20916 41636
rect 20860 41356 20916 41412
rect 21308 42530 21364 42532
rect 21308 42478 21310 42530
rect 21310 42478 21362 42530
rect 21362 42478 21364 42530
rect 21308 42476 21364 42478
rect 21532 41858 21588 41860
rect 21532 41806 21534 41858
rect 21534 41806 21586 41858
rect 21586 41806 21588 41858
rect 21532 41804 21588 41806
rect 22092 44546 22148 44548
rect 22092 44494 22094 44546
rect 22094 44494 22146 44546
rect 22146 44494 22148 44546
rect 22092 44492 22148 44494
rect 22316 43762 22372 43764
rect 22316 43710 22318 43762
rect 22318 43710 22370 43762
rect 22370 43710 22372 43762
rect 22316 43708 22372 43710
rect 21980 41916 22036 41972
rect 21980 41692 22036 41748
rect 21756 41410 21812 41412
rect 21756 41358 21758 41410
rect 21758 41358 21810 41410
rect 21810 41358 21812 41410
rect 21756 41356 21812 41358
rect 21420 41186 21476 41188
rect 21420 41134 21422 41186
rect 21422 41134 21474 41186
rect 21474 41134 21476 41186
rect 21420 41132 21476 41134
rect 21084 40626 21140 40628
rect 21084 40574 21086 40626
rect 21086 40574 21138 40626
rect 21138 40574 21140 40626
rect 21084 40572 21140 40574
rect 20636 40124 20692 40180
rect 21308 39788 21364 39844
rect 21980 41468 22036 41524
rect 22652 46172 22708 46228
rect 22764 45500 22820 45556
rect 23436 48188 23492 48244
rect 23436 47964 23492 48020
rect 23996 48188 24052 48244
rect 25228 49922 25284 49924
rect 25228 49870 25230 49922
rect 25230 49870 25282 49922
rect 25282 49870 25284 49922
rect 25228 49868 25284 49870
rect 24668 49026 24724 49028
rect 24668 48974 24670 49026
rect 24670 48974 24722 49026
rect 24722 48974 24724 49026
rect 24668 48972 24724 48974
rect 25564 49026 25620 49028
rect 25564 48974 25566 49026
rect 25566 48974 25618 49026
rect 25618 48974 25620 49026
rect 25564 48972 25620 48974
rect 25788 48300 25844 48356
rect 24556 48242 24612 48244
rect 24556 48190 24558 48242
rect 24558 48190 24610 48242
rect 24610 48190 24612 48242
rect 24556 48188 24612 48190
rect 24108 47628 24164 47684
rect 24668 47234 24724 47236
rect 24668 47182 24670 47234
rect 24670 47182 24722 47234
rect 24722 47182 24724 47234
rect 24668 47180 24724 47182
rect 25228 47180 25284 47236
rect 23996 46844 24052 46900
rect 24892 46844 24948 46900
rect 23660 46060 23716 46116
rect 23100 45388 23156 45444
rect 23436 45330 23492 45332
rect 23436 45278 23438 45330
rect 23438 45278 23490 45330
rect 23490 45278 23492 45330
rect 23436 45276 23492 45278
rect 23660 45164 23716 45220
rect 22988 44604 23044 44660
rect 22652 44210 22708 44212
rect 22652 44158 22654 44210
rect 22654 44158 22706 44210
rect 22706 44158 22708 44210
rect 22652 44156 22708 44158
rect 23100 44044 23156 44100
rect 23100 43426 23156 43428
rect 23100 43374 23102 43426
rect 23102 43374 23154 43426
rect 23154 43374 23156 43426
rect 23100 43372 23156 43374
rect 23212 42812 23268 42868
rect 22204 41804 22260 41860
rect 20860 38780 20916 38836
rect 19852 36594 19908 36596
rect 19852 36542 19854 36594
rect 19854 36542 19906 36594
rect 19906 36542 19908 36594
rect 19852 36540 19908 36542
rect 20412 36876 20468 36932
rect 20300 36258 20356 36260
rect 20300 36206 20302 36258
rect 20302 36206 20354 36258
rect 20354 36206 20356 36258
rect 20300 36204 20356 36206
rect 19836 36090 19892 36092
rect 19836 36038 19838 36090
rect 19838 36038 19890 36090
rect 19890 36038 19892 36090
rect 19836 36036 19892 36038
rect 19940 36090 19996 36092
rect 19940 36038 19942 36090
rect 19942 36038 19994 36090
rect 19994 36038 19996 36090
rect 19940 36036 19996 36038
rect 20044 36090 20100 36092
rect 20044 36038 20046 36090
rect 20046 36038 20098 36090
rect 20098 36038 20100 36090
rect 20044 36036 20100 36038
rect 19852 35868 19908 35924
rect 19404 35084 19460 35140
rect 20076 35532 20132 35588
rect 19964 35308 20020 35364
rect 19292 34412 19348 34468
rect 19180 33964 19236 34020
rect 19292 34076 19348 34132
rect 19068 33516 19124 33572
rect 19180 33404 19236 33460
rect 18620 33068 18676 33124
rect 17724 31388 17780 31444
rect 17836 31612 17892 31668
rect 17612 31276 17668 31332
rect 17612 31106 17668 31108
rect 17612 31054 17614 31106
rect 17614 31054 17666 31106
rect 17666 31054 17668 31106
rect 17612 31052 17668 31054
rect 17836 30940 17892 30996
rect 17724 30210 17780 30212
rect 17724 30158 17726 30210
rect 17726 30158 17778 30210
rect 17778 30158 17780 30210
rect 17724 30156 17780 30158
rect 17500 28700 17556 28756
rect 17500 27804 17556 27860
rect 17612 27020 17668 27076
rect 17388 26124 17444 26180
rect 17612 26796 17668 26852
rect 18172 31500 18228 31556
rect 18060 31218 18116 31220
rect 18060 31166 18062 31218
rect 18062 31166 18114 31218
rect 18114 31166 18116 31218
rect 18060 31164 18116 31166
rect 17948 30492 18004 30548
rect 18172 29820 18228 29876
rect 18956 33122 19012 33124
rect 18956 33070 18958 33122
rect 18958 33070 19010 33122
rect 19010 33070 19012 33122
rect 18956 33068 19012 33070
rect 19292 33292 19348 33348
rect 18844 31948 18900 32004
rect 18508 31778 18564 31780
rect 18508 31726 18510 31778
rect 18510 31726 18562 31778
rect 18562 31726 18564 31778
rect 18508 31724 18564 31726
rect 18508 31388 18564 31444
rect 18956 31388 19012 31444
rect 18732 31218 18788 31220
rect 18732 31166 18734 31218
rect 18734 31166 18786 31218
rect 18786 31166 18788 31218
rect 18732 31164 18788 31166
rect 19068 31218 19124 31220
rect 19068 31166 19070 31218
rect 19070 31166 19122 31218
rect 19122 31166 19124 31218
rect 19068 31164 19124 31166
rect 19180 32060 19236 32116
rect 18844 31106 18900 31108
rect 18844 31054 18846 31106
rect 18846 31054 18898 31106
rect 18898 31054 18900 31106
rect 18844 31052 18900 31054
rect 18956 30994 19012 30996
rect 18956 30942 18958 30994
rect 18958 30942 19010 30994
rect 19010 30942 19012 30994
rect 18956 30940 19012 30942
rect 19292 31388 19348 31444
rect 18396 29820 18452 29876
rect 18956 29820 19012 29876
rect 19292 30828 19348 30884
rect 19068 29708 19124 29764
rect 19068 29148 19124 29204
rect 19292 30604 19348 30660
rect 20748 36876 20804 36932
rect 20860 36428 20916 36484
rect 20300 35308 20356 35364
rect 19740 34636 19796 34692
rect 21084 37548 21140 37604
rect 21196 37212 21252 37268
rect 21084 37100 21140 37156
rect 20972 35980 21028 36036
rect 20860 35922 20916 35924
rect 20860 35870 20862 35922
rect 20862 35870 20914 35922
rect 20914 35870 20916 35922
rect 20860 35868 20916 35870
rect 20860 35420 20916 35476
rect 19836 34522 19892 34524
rect 19836 34470 19838 34522
rect 19838 34470 19890 34522
rect 19890 34470 19892 34522
rect 19836 34468 19892 34470
rect 19940 34522 19996 34524
rect 19940 34470 19942 34522
rect 19942 34470 19994 34522
rect 19994 34470 19996 34522
rect 19940 34468 19996 34470
rect 20044 34522 20100 34524
rect 20044 34470 20046 34522
rect 20046 34470 20098 34522
rect 20098 34470 20100 34522
rect 20044 34468 20100 34470
rect 19516 34130 19572 34132
rect 19516 34078 19518 34130
rect 19518 34078 19570 34130
rect 19570 34078 19572 34130
rect 19516 34076 19572 34078
rect 19516 33122 19572 33124
rect 19516 33070 19518 33122
rect 19518 33070 19570 33122
rect 19570 33070 19572 33122
rect 19516 33068 19572 33070
rect 19964 33068 20020 33124
rect 19836 32954 19892 32956
rect 19836 32902 19838 32954
rect 19838 32902 19890 32954
rect 19890 32902 19892 32954
rect 19836 32900 19892 32902
rect 19940 32954 19996 32956
rect 19940 32902 19942 32954
rect 19942 32902 19994 32954
rect 19994 32902 19996 32954
rect 19940 32900 19996 32902
rect 20044 32954 20100 32956
rect 20044 32902 20046 32954
rect 20046 32902 20098 32954
rect 20098 32902 20100 32954
rect 20044 32900 20100 32902
rect 20300 33964 20356 34020
rect 20300 32956 20356 33012
rect 20188 32844 20244 32900
rect 19516 32620 19572 32676
rect 19852 32060 19908 32116
rect 19964 32396 20020 32452
rect 19516 31612 19572 31668
rect 20972 35308 21028 35364
rect 20972 34412 21028 34468
rect 20972 34130 21028 34132
rect 20972 34078 20974 34130
rect 20974 34078 21026 34130
rect 21026 34078 21028 34130
rect 20972 34076 21028 34078
rect 21532 38834 21588 38836
rect 21532 38782 21534 38834
rect 21534 38782 21586 38834
rect 21586 38782 21588 38834
rect 21532 38780 21588 38782
rect 21420 37436 21476 37492
rect 21420 37154 21476 37156
rect 21420 37102 21422 37154
rect 21422 37102 21474 37154
rect 21474 37102 21476 37154
rect 21420 37100 21476 37102
rect 21532 36988 21588 37044
rect 22540 41020 22596 41076
rect 21980 40572 22036 40628
rect 22316 40460 22372 40516
rect 22540 40402 22596 40404
rect 22540 40350 22542 40402
rect 22542 40350 22594 40402
rect 22594 40350 22596 40402
rect 22540 40348 22596 40350
rect 23100 42476 23156 42532
rect 22876 42140 22932 42196
rect 23436 44268 23492 44324
rect 24332 44994 24388 44996
rect 24332 44942 24334 44994
rect 24334 44942 24386 44994
rect 24386 44942 24388 44994
rect 24332 44940 24388 44942
rect 24332 44604 24388 44660
rect 23660 44156 23716 44212
rect 24220 44210 24276 44212
rect 24220 44158 24222 44210
rect 24222 44158 24274 44210
rect 24274 44158 24276 44210
rect 24220 44156 24276 44158
rect 23772 43820 23828 43876
rect 23548 43596 23604 43652
rect 23996 43596 24052 43652
rect 24220 43538 24276 43540
rect 24220 43486 24222 43538
rect 24222 43486 24274 43538
rect 24274 43486 24276 43538
rect 24220 43484 24276 43486
rect 24220 43260 24276 43316
rect 24108 43036 24164 43092
rect 23100 41356 23156 41412
rect 23212 41580 23268 41636
rect 23324 41804 23380 41860
rect 23324 41020 23380 41076
rect 23436 41692 23492 41748
rect 23212 40572 23268 40628
rect 23436 40348 23492 40404
rect 22652 40124 22708 40180
rect 22204 39788 22260 39844
rect 22092 38892 22148 38948
rect 21980 38834 22036 38836
rect 21980 38782 21982 38834
rect 21982 38782 22034 38834
rect 22034 38782 22036 38834
rect 21980 38780 22036 38782
rect 21980 38220 22036 38276
rect 21980 37548 22036 37604
rect 21980 37324 22036 37380
rect 21868 36540 21924 36596
rect 21420 35532 21476 35588
rect 21644 35532 21700 35588
rect 21308 34076 21364 34132
rect 21196 33740 21252 33796
rect 20636 33180 20692 33236
rect 20076 31836 20132 31892
rect 20188 31778 20244 31780
rect 20188 31726 20190 31778
rect 20190 31726 20242 31778
rect 20242 31726 20244 31778
rect 20188 31724 20244 31726
rect 18620 28924 18676 28980
rect 18172 28364 18228 28420
rect 20300 31554 20356 31556
rect 20300 31502 20302 31554
rect 20302 31502 20354 31554
rect 20354 31502 20356 31554
rect 20300 31500 20356 31502
rect 19836 31386 19892 31388
rect 19836 31334 19838 31386
rect 19838 31334 19890 31386
rect 19890 31334 19892 31386
rect 19836 31332 19892 31334
rect 19940 31386 19996 31388
rect 19940 31334 19942 31386
rect 19942 31334 19994 31386
rect 19994 31334 19996 31386
rect 19940 31332 19996 31334
rect 20044 31386 20100 31388
rect 20044 31334 20046 31386
rect 20046 31334 20098 31386
rect 20098 31334 20100 31386
rect 20044 31332 20100 31334
rect 20860 33628 20916 33684
rect 21868 34524 21924 34580
rect 22652 38668 22708 38724
rect 22540 37212 22596 37268
rect 22876 38332 22932 38388
rect 22876 38162 22932 38164
rect 22876 38110 22878 38162
rect 22878 38110 22930 38162
rect 22930 38110 22932 38162
rect 22876 38108 22932 38110
rect 22764 37548 22820 37604
rect 22764 37324 22820 37380
rect 22988 36988 23044 37044
rect 22540 36092 22596 36148
rect 22876 35868 22932 35924
rect 21868 34076 21924 34132
rect 21644 33628 21700 33684
rect 20860 33068 20916 33124
rect 21644 32732 21700 32788
rect 20860 32620 20916 32676
rect 19740 31164 19796 31220
rect 18732 28812 18788 28868
rect 18844 28588 18900 28644
rect 17836 27804 17892 27860
rect 18060 27356 18116 27412
rect 18396 27580 18452 27636
rect 18508 27804 18564 27860
rect 17948 27186 18004 27188
rect 17948 27134 17950 27186
rect 17950 27134 18002 27186
rect 18002 27134 18004 27186
rect 17948 27132 18004 27134
rect 18172 27020 18228 27076
rect 17948 26572 18004 26628
rect 17612 26402 17668 26404
rect 17612 26350 17614 26402
rect 17614 26350 17666 26402
rect 17666 26350 17668 26402
rect 17612 26348 17668 26350
rect 17948 26290 18004 26292
rect 17948 26238 17950 26290
rect 17950 26238 18002 26290
rect 18002 26238 18004 26290
rect 17948 26236 18004 26238
rect 17388 25116 17444 25172
rect 17612 25788 17668 25844
rect 17276 24892 17332 24948
rect 17724 25228 17780 25284
rect 17836 24722 17892 24724
rect 17836 24670 17838 24722
rect 17838 24670 17890 24722
rect 17890 24670 17892 24722
rect 17836 24668 17892 24670
rect 16828 24556 16884 24612
rect 18732 27132 18788 27188
rect 19180 28754 19236 28756
rect 19180 28702 19182 28754
rect 19182 28702 19234 28754
rect 19234 28702 19236 28754
rect 19180 28700 19236 28702
rect 19068 27580 19124 27636
rect 20636 31500 20692 31556
rect 20076 30716 20132 30772
rect 19964 30380 20020 30436
rect 19964 30098 20020 30100
rect 19964 30046 19966 30098
rect 19966 30046 20018 30098
rect 20018 30046 20020 30098
rect 19964 30044 20020 30046
rect 20076 29932 20132 29988
rect 19836 29818 19892 29820
rect 19836 29766 19838 29818
rect 19838 29766 19890 29818
rect 19890 29766 19892 29818
rect 19836 29764 19892 29766
rect 19940 29818 19996 29820
rect 19940 29766 19942 29818
rect 19942 29766 19994 29818
rect 19994 29766 19996 29818
rect 19940 29764 19996 29766
rect 20044 29818 20100 29820
rect 20044 29766 20046 29818
rect 20046 29766 20098 29818
rect 20098 29766 20100 29818
rect 20044 29764 20100 29766
rect 19740 29596 19796 29652
rect 19292 27916 19348 27972
rect 19404 27858 19460 27860
rect 19404 27806 19406 27858
rect 19406 27806 19458 27858
rect 19458 27806 19460 27858
rect 19404 27804 19460 27806
rect 20076 29650 20132 29652
rect 20076 29598 20078 29650
rect 20078 29598 20130 29650
rect 20130 29598 20132 29650
rect 20076 29596 20132 29598
rect 21420 32450 21476 32452
rect 21420 32398 21422 32450
rect 21422 32398 21474 32450
rect 21474 32398 21476 32450
rect 21420 32396 21476 32398
rect 21084 32284 21140 32340
rect 20860 31890 20916 31892
rect 20860 31838 20862 31890
rect 20862 31838 20914 31890
rect 20914 31838 20916 31890
rect 20860 31836 20916 31838
rect 20412 29538 20468 29540
rect 20412 29486 20414 29538
rect 20414 29486 20466 29538
rect 20466 29486 20468 29538
rect 20412 29484 20468 29486
rect 20748 30156 20804 30212
rect 19964 28924 20020 28980
rect 20076 29148 20132 29204
rect 20188 29036 20244 29092
rect 20188 28364 20244 28420
rect 19836 28250 19892 28252
rect 19836 28198 19838 28250
rect 19838 28198 19890 28250
rect 19890 28198 19892 28250
rect 19836 28196 19892 28198
rect 19940 28250 19996 28252
rect 19940 28198 19942 28250
rect 19942 28198 19994 28250
rect 19994 28198 19996 28250
rect 19940 28196 19996 28198
rect 20044 28250 20100 28252
rect 20044 28198 20046 28250
rect 20046 28198 20098 28250
rect 20098 28198 20100 28250
rect 20044 28196 20100 28198
rect 19964 27858 20020 27860
rect 19964 27806 19966 27858
rect 19966 27806 20018 27858
rect 20018 27806 20020 27858
rect 19964 27804 20020 27806
rect 20524 27970 20580 27972
rect 20524 27918 20526 27970
rect 20526 27918 20578 27970
rect 20578 27918 20580 27970
rect 20524 27916 20580 27918
rect 20972 30268 21028 30324
rect 21420 31666 21476 31668
rect 21420 31614 21422 31666
rect 21422 31614 21474 31666
rect 21474 31614 21476 31666
rect 21420 31612 21476 31614
rect 21420 31276 21476 31332
rect 21420 30716 21476 30772
rect 21420 30434 21476 30436
rect 21420 30382 21422 30434
rect 21422 30382 21474 30434
rect 21474 30382 21476 30434
rect 21420 30380 21476 30382
rect 21868 31724 21924 31780
rect 22764 34748 22820 34804
rect 22652 34636 22708 34692
rect 22876 35308 22932 35364
rect 22092 33404 22148 33460
rect 22652 33852 22708 33908
rect 22092 33180 22148 33236
rect 22092 32172 22148 32228
rect 21868 31500 21924 31556
rect 21196 29708 21252 29764
rect 21308 29596 21364 29652
rect 21084 29484 21140 29540
rect 20972 29426 21028 29428
rect 20972 29374 20974 29426
rect 20974 29374 21026 29426
rect 21026 29374 21028 29426
rect 20972 29372 21028 29374
rect 20188 27468 20244 27524
rect 18284 26962 18340 26964
rect 18284 26910 18286 26962
rect 18286 26910 18338 26962
rect 18338 26910 18340 26962
rect 18284 26908 18340 26910
rect 18508 26402 18564 26404
rect 18508 26350 18510 26402
rect 18510 26350 18562 26402
rect 18562 26350 18564 26402
rect 18508 26348 18564 26350
rect 18172 23826 18228 23828
rect 18172 23774 18174 23826
rect 18174 23774 18226 23826
rect 18226 23774 18228 23826
rect 18172 23772 18228 23774
rect 18844 25506 18900 25508
rect 18844 25454 18846 25506
rect 18846 25454 18898 25506
rect 18898 25454 18900 25506
rect 18844 25452 18900 25454
rect 18620 25282 18676 25284
rect 18620 25230 18622 25282
rect 18622 25230 18674 25282
rect 18674 25230 18676 25282
rect 18620 25228 18676 25230
rect 20300 26796 20356 26852
rect 19836 26682 19892 26684
rect 19836 26630 19838 26682
rect 19838 26630 19890 26682
rect 19890 26630 19892 26682
rect 19836 26628 19892 26630
rect 19940 26682 19996 26684
rect 19940 26630 19942 26682
rect 19942 26630 19994 26682
rect 19994 26630 19996 26682
rect 19940 26628 19996 26630
rect 20044 26682 20100 26684
rect 20044 26630 20046 26682
rect 20046 26630 20098 26682
rect 20098 26630 20100 26682
rect 20044 26628 20100 26630
rect 19180 26124 19236 26180
rect 19852 26178 19908 26180
rect 19852 26126 19854 26178
rect 19854 26126 19906 26178
rect 19906 26126 19908 26178
rect 19852 26124 19908 26126
rect 19740 25564 19796 25620
rect 19964 25788 20020 25844
rect 20300 25564 20356 25620
rect 19852 25452 19908 25508
rect 19068 25228 19124 25284
rect 20076 25228 20132 25284
rect 19836 25114 19892 25116
rect 19836 25062 19838 25114
rect 19838 25062 19890 25114
rect 19890 25062 19892 25114
rect 19836 25060 19892 25062
rect 19940 25114 19996 25116
rect 19940 25062 19942 25114
rect 19942 25062 19994 25114
rect 19994 25062 19996 25114
rect 19940 25060 19996 25062
rect 20044 25114 20100 25116
rect 20044 25062 20046 25114
rect 20046 25062 20098 25114
rect 20098 25062 20100 25114
rect 20044 25060 20100 25062
rect 18508 24610 18564 24612
rect 18508 24558 18510 24610
rect 18510 24558 18562 24610
rect 18562 24558 18564 24610
rect 18508 24556 18564 24558
rect 19068 24556 19124 24612
rect 16156 22876 16212 22932
rect 17612 22876 17668 22932
rect 19964 24668 20020 24724
rect 19740 24050 19796 24052
rect 19740 23998 19742 24050
rect 19742 23998 19794 24050
rect 19794 23998 19796 24050
rect 19740 23996 19796 23998
rect 20188 23938 20244 23940
rect 20188 23886 20190 23938
rect 20190 23886 20242 23938
rect 20242 23886 20244 23938
rect 20188 23884 20244 23886
rect 20748 26178 20804 26180
rect 20748 26126 20750 26178
rect 20750 26126 20802 26178
rect 20802 26126 20804 26178
rect 20748 26124 20804 26126
rect 21532 29426 21588 29428
rect 21532 29374 21534 29426
rect 21534 29374 21586 29426
rect 21586 29374 21588 29426
rect 21532 29372 21588 29374
rect 21980 29596 22036 29652
rect 21980 29426 22036 29428
rect 21980 29374 21982 29426
rect 21982 29374 22034 29426
rect 22034 29374 22036 29426
rect 21980 29372 22036 29374
rect 21532 28530 21588 28532
rect 21532 28478 21534 28530
rect 21534 28478 21586 28530
rect 21586 28478 21588 28530
rect 21532 28476 21588 28478
rect 21084 26460 21140 26516
rect 21644 27970 21700 27972
rect 21644 27918 21646 27970
rect 21646 27918 21698 27970
rect 21698 27918 21700 27970
rect 21644 27916 21700 27918
rect 21420 26908 21476 26964
rect 20524 23996 20580 24052
rect 21084 23884 21140 23940
rect 19836 23546 19892 23548
rect 19836 23494 19838 23546
rect 19838 23494 19890 23546
rect 19890 23494 19892 23546
rect 19836 23492 19892 23494
rect 19940 23546 19996 23548
rect 19940 23494 19942 23546
rect 19942 23494 19994 23546
rect 19994 23494 19996 23546
rect 19940 23492 19996 23494
rect 20044 23546 20100 23548
rect 20044 23494 20046 23546
rect 20046 23494 20098 23546
rect 20098 23494 20100 23546
rect 20044 23492 20100 23494
rect 21084 23548 21140 23604
rect 21644 26290 21700 26292
rect 21644 26238 21646 26290
rect 21646 26238 21698 26290
rect 21698 26238 21700 26290
rect 21644 26236 21700 26238
rect 22092 26290 22148 26292
rect 22092 26238 22094 26290
rect 22094 26238 22146 26290
rect 22146 26238 22148 26290
rect 22092 26236 22148 26238
rect 21532 25282 21588 25284
rect 21532 25230 21534 25282
rect 21534 25230 21586 25282
rect 21586 25230 21588 25282
rect 21532 25228 21588 25230
rect 22092 24834 22148 24836
rect 22092 24782 22094 24834
rect 22094 24782 22146 24834
rect 22146 24782 22148 24834
rect 22092 24780 22148 24782
rect 22316 33292 22372 33348
rect 22540 32508 22596 32564
rect 22316 31778 22372 31780
rect 22316 31726 22318 31778
rect 22318 31726 22370 31778
rect 22370 31726 22372 31778
rect 22316 31724 22372 31726
rect 22540 31724 22596 31780
rect 22764 32956 22820 33012
rect 22764 31778 22820 31780
rect 22764 31726 22766 31778
rect 22766 31726 22818 31778
rect 22818 31726 22820 31778
rect 22764 31724 22820 31726
rect 22988 33404 23044 33460
rect 23212 38722 23268 38724
rect 23212 38670 23214 38722
rect 23214 38670 23266 38722
rect 23266 38670 23268 38722
rect 23212 38668 23268 38670
rect 23324 38556 23380 38612
rect 23324 37996 23380 38052
rect 23660 42476 23716 42532
rect 23996 42530 24052 42532
rect 23996 42478 23998 42530
rect 23998 42478 24050 42530
rect 24050 42478 24052 42530
rect 23996 42476 24052 42478
rect 23884 42364 23940 42420
rect 23660 42252 23716 42308
rect 23884 40460 23940 40516
rect 23884 39506 23940 39508
rect 23884 39454 23886 39506
rect 23886 39454 23938 39506
rect 23938 39454 23940 39506
rect 23884 39452 23940 39454
rect 24220 42252 24276 42308
rect 24556 45778 24612 45780
rect 24556 45726 24558 45778
rect 24558 45726 24610 45778
rect 24610 45726 24612 45778
rect 24556 45724 24612 45726
rect 24668 45164 24724 45220
rect 24668 44604 24724 44660
rect 24668 44434 24724 44436
rect 24668 44382 24670 44434
rect 24670 44382 24722 44434
rect 24722 44382 24724 44434
rect 24668 44380 24724 44382
rect 24556 44268 24612 44324
rect 24556 43820 24612 43876
rect 24668 43314 24724 43316
rect 24668 43262 24670 43314
rect 24670 43262 24722 43314
rect 24722 43262 24724 43314
rect 24668 43260 24724 43262
rect 25004 44098 25060 44100
rect 25004 44046 25006 44098
rect 25006 44046 25058 44098
rect 25058 44046 25060 44098
rect 25004 44044 25060 44046
rect 24444 42754 24500 42756
rect 24444 42702 24446 42754
rect 24446 42702 24498 42754
rect 24498 42702 24500 42754
rect 24444 42700 24500 42702
rect 24668 42364 24724 42420
rect 25004 42700 25060 42756
rect 24668 41468 24724 41524
rect 24892 41356 24948 41412
rect 24668 39340 24724 39396
rect 24220 38946 24276 38948
rect 24220 38894 24222 38946
rect 24222 38894 24274 38946
rect 24274 38894 24276 38946
rect 24220 38892 24276 38894
rect 24108 38220 24164 38276
rect 23212 36876 23268 36932
rect 23436 36876 23492 36932
rect 23548 35868 23604 35924
rect 23324 33458 23380 33460
rect 23324 33406 23326 33458
rect 23326 33406 23378 33458
rect 23378 33406 23380 33458
rect 23324 33404 23380 33406
rect 23772 35196 23828 35252
rect 23884 35308 23940 35364
rect 23772 34524 23828 34580
rect 24332 37884 24388 37940
rect 24108 37772 24164 37828
rect 24220 36316 24276 36372
rect 24108 34972 24164 35028
rect 23772 33852 23828 33908
rect 23436 33292 23492 33348
rect 23212 33122 23268 33124
rect 23212 33070 23214 33122
rect 23214 33070 23266 33122
rect 23266 33070 23268 33122
rect 23212 33068 23268 33070
rect 23436 32732 23492 32788
rect 23100 32620 23156 32676
rect 22988 32508 23044 32564
rect 22988 31836 23044 31892
rect 23436 32172 23492 32228
rect 22652 31276 22708 31332
rect 22540 30044 22596 30100
rect 22652 29820 22708 29876
rect 22428 29538 22484 29540
rect 22428 29486 22430 29538
rect 22430 29486 22482 29538
rect 22482 29486 22484 29538
rect 22428 29484 22484 29486
rect 22876 28476 22932 28532
rect 22652 27746 22708 27748
rect 22652 27694 22654 27746
rect 22654 27694 22706 27746
rect 22706 27694 22708 27746
rect 22652 27692 22708 27694
rect 23100 31612 23156 31668
rect 23996 34130 24052 34132
rect 23996 34078 23998 34130
rect 23998 34078 24050 34130
rect 24050 34078 24052 34130
rect 23996 34076 24052 34078
rect 23660 31724 23716 31780
rect 23212 31276 23268 31332
rect 23212 30828 23268 30884
rect 23212 30098 23268 30100
rect 23212 30046 23214 30098
rect 23214 30046 23266 30098
rect 23266 30046 23268 30098
rect 23212 30044 23268 30046
rect 23100 29372 23156 29428
rect 24332 35756 24388 35812
rect 24220 32956 24276 33012
rect 24444 32956 24500 33012
rect 24556 37548 24612 37604
rect 24332 31948 24388 32004
rect 23884 31218 23940 31220
rect 23884 31166 23886 31218
rect 23886 31166 23938 31218
rect 23938 31166 23940 31218
rect 23884 31164 23940 31166
rect 24220 30994 24276 30996
rect 24220 30942 24222 30994
rect 24222 30942 24274 30994
rect 24274 30942 24276 30994
rect 24220 30940 24276 30942
rect 23548 30210 23604 30212
rect 23548 30158 23550 30210
rect 23550 30158 23602 30210
rect 23602 30158 23604 30210
rect 23548 30156 23604 30158
rect 23548 29932 23604 29988
rect 23436 29820 23492 29876
rect 23436 28588 23492 28644
rect 23548 27692 23604 27748
rect 24444 31724 24500 31780
rect 24444 31500 24500 31556
rect 24444 31106 24500 31108
rect 24444 31054 24446 31106
rect 24446 31054 24498 31106
rect 24498 31054 24500 31106
rect 24444 31052 24500 31054
rect 24668 37324 24724 37380
rect 24668 34972 24724 35028
rect 24668 32450 24724 32452
rect 24668 32398 24670 32450
rect 24670 32398 24722 32450
rect 24722 32398 24724 32450
rect 24668 32396 24724 32398
rect 24108 30098 24164 30100
rect 24108 30046 24110 30098
rect 24110 30046 24162 30098
rect 24162 30046 24164 30098
rect 24108 30044 24164 30046
rect 23884 29708 23940 29764
rect 23772 27186 23828 27188
rect 23772 27134 23774 27186
rect 23774 27134 23826 27186
rect 23826 27134 23828 27186
rect 23772 27132 23828 27134
rect 22204 24668 22260 24724
rect 21868 23548 21924 23604
rect 23100 26236 23156 26292
rect 22652 25340 22708 25396
rect 22764 25676 22820 25732
rect 22540 25228 22596 25284
rect 23100 25116 23156 25172
rect 23324 25788 23380 25844
rect 22316 24108 22372 24164
rect 23548 25676 23604 25732
rect 23660 25506 23716 25508
rect 23660 25454 23662 25506
rect 23662 25454 23714 25506
rect 23714 25454 23716 25506
rect 23660 25452 23716 25454
rect 23548 25394 23604 25396
rect 23548 25342 23550 25394
rect 23550 25342 23602 25394
rect 23602 25342 23604 25394
rect 23548 25340 23604 25342
rect 23772 24220 23828 24276
rect 24108 29650 24164 29652
rect 24108 29598 24110 29650
rect 24110 29598 24162 29650
rect 24162 29598 24164 29650
rect 24108 29596 24164 29598
rect 24556 30156 24612 30212
rect 24332 29708 24388 29764
rect 24444 29260 24500 29316
rect 24220 28530 24276 28532
rect 24220 28478 24222 28530
rect 24222 28478 24274 28530
rect 24274 28478 24276 28530
rect 24220 28476 24276 28478
rect 24332 28418 24388 28420
rect 24332 28366 24334 28418
rect 24334 28366 24386 28418
rect 24386 28366 24388 28418
rect 24332 28364 24388 28366
rect 24668 28028 24724 28084
rect 24668 27580 24724 27636
rect 25564 44940 25620 44996
rect 26012 48300 26068 48356
rect 27580 51212 27636 51268
rect 27356 50706 27412 50708
rect 27356 50654 27358 50706
rect 27358 50654 27410 50706
rect 27410 50654 27412 50706
rect 27356 50652 27412 50654
rect 29372 52162 29428 52164
rect 29372 52110 29374 52162
rect 29374 52110 29426 52162
rect 29426 52110 29428 52162
rect 29372 52108 29428 52110
rect 28252 51266 28308 51268
rect 28252 51214 28254 51266
rect 28254 51214 28306 51266
rect 28306 51214 28308 51266
rect 28252 51212 28308 51214
rect 27132 48860 27188 48916
rect 26572 48242 26628 48244
rect 26572 48190 26574 48242
rect 26574 48190 26626 48242
rect 26626 48190 26628 48242
rect 26572 48188 26628 48190
rect 25900 45218 25956 45220
rect 25900 45166 25902 45218
rect 25902 45166 25954 45218
rect 25954 45166 25956 45218
rect 25900 45164 25956 45166
rect 26796 45890 26852 45892
rect 26796 45838 26798 45890
rect 26798 45838 26850 45890
rect 26850 45838 26852 45890
rect 26796 45836 26852 45838
rect 26124 45106 26180 45108
rect 26124 45054 26126 45106
rect 26126 45054 26178 45106
rect 26178 45054 26180 45106
rect 26124 45052 26180 45054
rect 26124 44434 26180 44436
rect 26124 44382 26126 44434
rect 26126 44382 26178 44434
rect 26178 44382 26180 44434
rect 26124 44380 26180 44382
rect 25564 43372 25620 43428
rect 25564 42754 25620 42756
rect 25564 42702 25566 42754
rect 25566 42702 25618 42754
rect 25618 42702 25620 42754
rect 25564 42700 25620 42702
rect 25452 42642 25508 42644
rect 25452 42590 25454 42642
rect 25454 42590 25506 42642
rect 25506 42590 25508 42642
rect 25452 42588 25508 42590
rect 26348 44604 26404 44660
rect 27132 45500 27188 45556
rect 27020 44380 27076 44436
rect 26684 44322 26740 44324
rect 26684 44270 26686 44322
rect 26686 44270 26738 44322
rect 26738 44270 26740 44322
rect 26684 44268 26740 44270
rect 26460 44210 26516 44212
rect 26460 44158 26462 44210
rect 26462 44158 26514 44210
rect 26514 44158 26516 44210
rect 26460 44156 26516 44158
rect 25452 42364 25508 42420
rect 25116 40572 25172 40628
rect 25340 41692 25396 41748
rect 25004 39228 25060 39284
rect 25116 39058 25172 39060
rect 25116 39006 25118 39058
rect 25118 39006 25170 39058
rect 25170 39006 25172 39058
rect 25116 39004 25172 39006
rect 25340 39228 25396 39284
rect 25564 39228 25620 39284
rect 25676 40178 25732 40180
rect 25676 40126 25678 40178
rect 25678 40126 25730 40178
rect 25730 40126 25732 40178
rect 25676 40124 25732 40126
rect 24892 37884 24948 37940
rect 25004 38444 25060 38500
rect 25228 37490 25284 37492
rect 25228 37438 25230 37490
rect 25230 37438 25282 37490
rect 25282 37438 25284 37490
rect 25228 37436 25284 37438
rect 25228 37100 25284 37156
rect 25564 38722 25620 38724
rect 25564 38670 25566 38722
rect 25566 38670 25618 38722
rect 25618 38670 25620 38722
rect 25564 38668 25620 38670
rect 25564 38108 25620 38164
rect 25452 37212 25508 37268
rect 25788 39340 25844 39396
rect 26348 43932 26404 43988
rect 26572 43650 26628 43652
rect 26572 43598 26574 43650
rect 26574 43598 26626 43650
rect 26626 43598 26628 43650
rect 26572 43596 26628 43598
rect 26796 42476 26852 42532
rect 26572 41858 26628 41860
rect 26572 41806 26574 41858
rect 26574 41806 26626 41858
rect 26626 41806 26628 41858
rect 26572 41804 26628 41806
rect 26348 40460 26404 40516
rect 26460 41020 26516 41076
rect 26348 40178 26404 40180
rect 26348 40126 26350 40178
rect 26350 40126 26402 40178
rect 26402 40126 26404 40178
rect 26348 40124 26404 40126
rect 25900 39004 25956 39060
rect 26124 40012 26180 40068
rect 27356 47458 27412 47460
rect 27356 47406 27358 47458
rect 27358 47406 27410 47458
rect 27410 47406 27412 47458
rect 27356 47404 27412 47406
rect 27356 45778 27412 45780
rect 27356 45726 27358 45778
rect 27358 45726 27410 45778
rect 27410 45726 27412 45778
rect 27356 45724 27412 45726
rect 27692 47404 27748 47460
rect 29596 51996 29652 52052
rect 33180 55298 33236 55300
rect 33180 55246 33182 55298
rect 33182 55246 33234 55298
rect 33234 55246 33236 55298
rect 33180 55244 33236 55246
rect 33628 55298 33684 55300
rect 33628 55246 33630 55298
rect 33630 55246 33682 55298
rect 33682 55246 33684 55298
rect 33628 55244 33684 55246
rect 32508 54402 32564 54404
rect 32508 54350 32510 54402
rect 32510 54350 32562 54402
rect 32562 54350 32564 54402
rect 32508 54348 32564 54350
rect 32060 53676 32116 53732
rect 32284 53058 32340 53060
rect 32284 53006 32286 53058
rect 32286 53006 32338 53058
rect 32338 53006 32340 53058
rect 32284 53004 32340 53006
rect 30828 52780 30884 52836
rect 31948 52834 32004 52836
rect 31948 52782 31950 52834
rect 31950 52782 32002 52834
rect 32002 52782 32004 52834
rect 31948 52780 32004 52782
rect 30492 51324 30548 51380
rect 32620 53618 32676 53620
rect 32620 53566 32622 53618
rect 32622 53566 32674 53618
rect 32674 53566 32676 53618
rect 32620 53564 32676 53566
rect 33068 53564 33124 53620
rect 33404 54348 33460 54404
rect 33292 53788 33348 53844
rect 33180 52946 33236 52948
rect 33180 52894 33182 52946
rect 33182 52894 33234 52946
rect 33234 52894 33236 52946
rect 33180 52892 33236 52894
rect 32844 52274 32900 52276
rect 32844 52222 32846 52274
rect 32846 52222 32898 52274
rect 32898 52222 32900 52274
rect 32844 52220 32900 52222
rect 32508 51324 32564 51380
rect 30380 51100 30436 51156
rect 30380 49980 30436 50036
rect 29260 49756 29316 49812
rect 29260 49084 29316 49140
rect 29484 48354 29540 48356
rect 29484 48302 29486 48354
rect 29486 48302 29538 48354
rect 29538 48302 29540 48354
rect 29484 48300 29540 48302
rect 29036 48242 29092 48244
rect 29036 48190 29038 48242
rect 29038 48190 29090 48242
rect 29090 48190 29092 48242
rect 29036 48188 29092 48190
rect 28588 48076 28644 48132
rect 29484 47964 29540 48020
rect 27916 46956 27972 47012
rect 28812 46732 28868 46788
rect 28140 45500 28196 45556
rect 28252 46060 28308 46116
rect 27468 44098 27524 44100
rect 27468 44046 27470 44098
rect 27470 44046 27522 44098
rect 27522 44046 27524 44098
rect 27468 44044 27524 44046
rect 28364 45612 28420 45668
rect 26908 41804 26964 41860
rect 27356 42028 27412 42084
rect 27020 41132 27076 41188
rect 27132 41692 27188 41748
rect 27132 40796 27188 40852
rect 27356 40908 27412 40964
rect 27356 40626 27412 40628
rect 27356 40574 27358 40626
rect 27358 40574 27410 40626
rect 27410 40574 27412 40626
rect 27356 40572 27412 40574
rect 27244 40460 27300 40516
rect 26572 40348 26628 40404
rect 26124 39564 26180 39620
rect 25788 38668 25844 38724
rect 26348 39228 26404 39284
rect 25676 37548 25732 37604
rect 26236 38722 26292 38724
rect 26236 38670 26238 38722
rect 26238 38670 26290 38722
rect 26290 38670 26292 38722
rect 26236 38668 26292 38670
rect 26236 38162 26292 38164
rect 26236 38110 26238 38162
rect 26238 38110 26290 38162
rect 26290 38110 26292 38162
rect 26236 38108 26292 38110
rect 26012 37996 26068 38052
rect 25564 37100 25620 37156
rect 25340 36652 25396 36708
rect 25788 36988 25844 37044
rect 25340 36482 25396 36484
rect 25340 36430 25342 36482
rect 25342 36430 25394 36482
rect 25394 36430 25396 36482
rect 25340 36428 25396 36430
rect 26236 37378 26292 37380
rect 26236 37326 26238 37378
rect 26238 37326 26290 37378
rect 26290 37326 26292 37378
rect 26236 37324 26292 37326
rect 26124 36876 26180 36932
rect 26012 36652 26068 36708
rect 25676 35868 25732 35924
rect 25340 35756 25396 35812
rect 25340 35196 25396 35252
rect 25452 34860 25508 34916
rect 25228 33404 25284 33460
rect 25340 33628 25396 33684
rect 25116 33292 25172 33348
rect 25340 33180 25396 33236
rect 25340 32562 25396 32564
rect 25340 32510 25342 32562
rect 25342 32510 25394 32562
rect 25394 32510 25396 32562
rect 25340 32508 25396 32510
rect 25564 32396 25620 32452
rect 26012 35308 26068 35364
rect 26236 35196 26292 35252
rect 26684 39564 26740 39620
rect 27132 39506 27188 39508
rect 27132 39454 27134 39506
rect 27134 39454 27186 39506
rect 27186 39454 27188 39506
rect 27132 39452 27188 39454
rect 27020 39340 27076 39396
rect 26684 39228 26740 39284
rect 27132 38892 27188 38948
rect 26908 38834 26964 38836
rect 26908 38782 26910 38834
rect 26910 38782 26962 38834
rect 26962 38782 26964 38834
rect 26908 38780 26964 38782
rect 28252 42700 28308 42756
rect 28700 45218 28756 45220
rect 28700 45166 28702 45218
rect 28702 45166 28754 45218
rect 28754 45166 28756 45218
rect 28700 45164 28756 45166
rect 28476 44156 28532 44212
rect 28588 43148 28644 43204
rect 27916 42588 27972 42644
rect 27804 41692 27860 41748
rect 28364 41692 28420 41748
rect 27916 41298 27972 41300
rect 27916 41246 27918 41298
rect 27918 41246 27970 41298
rect 27970 41246 27972 41298
rect 27916 41244 27972 41246
rect 27692 40796 27748 40852
rect 27580 40684 27636 40740
rect 27804 40460 27860 40516
rect 28364 40348 28420 40404
rect 28476 41132 28532 41188
rect 27916 40236 27972 40292
rect 28252 40124 28308 40180
rect 28028 39900 28084 39956
rect 27916 38946 27972 38948
rect 27916 38894 27918 38946
rect 27918 38894 27970 38946
rect 27970 38894 27972 38946
rect 27916 38892 27972 38894
rect 27692 38668 27748 38724
rect 28252 39564 28308 39620
rect 28588 40684 28644 40740
rect 29148 43932 29204 43988
rect 29260 46284 29316 46340
rect 29148 43650 29204 43652
rect 29148 43598 29150 43650
rect 29150 43598 29202 43650
rect 29202 43598 29204 43650
rect 29148 43596 29204 43598
rect 29148 40908 29204 40964
rect 26572 38220 26628 38276
rect 27244 38332 27300 38388
rect 26796 37490 26852 37492
rect 26796 37438 26798 37490
rect 26798 37438 26850 37490
rect 26850 37438 26852 37490
rect 26796 37436 26852 37438
rect 26572 37266 26628 37268
rect 26572 37214 26574 37266
rect 26574 37214 26626 37266
rect 26626 37214 26628 37266
rect 26572 37212 26628 37214
rect 27692 37772 27748 37828
rect 27468 37212 27524 37268
rect 26572 36764 26628 36820
rect 26460 35026 26516 35028
rect 26460 34974 26462 35026
rect 26462 34974 26514 35026
rect 26514 34974 26516 35026
rect 26460 34972 26516 34974
rect 26236 34188 26292 34244
rect 26460 33852 26516 33908
rect 26684 35420 26740 35476
rect 26908 36876 26964 36932
rect 26684 34914 26740 34916
rect 26684 34862 26686 34914
rect 26686 34862 26738 34914
rect 26738 34862 26740 34914
rect 26684 34860 26740 34862
rect 26796 34076 26852 34132
rect 26572 32620 26628 32676
rect 26124 31276 26180 31332
rect 26348 31218 26404 31220
rect 26348 31166 26350 31218
rect 26350 31166 26402 31218
rect 26402 31166 26404 31218
rect 26348 31164 26404 31166
rect 25676 30604 25732 30660
rect 25228 30210 25284 30212
rect 25228 30158 25230 30210
rect 25230 30158 25282 30210
rect 25282 30158 25284 30210
rect 25228 30156 25284 30158
rect 25116 30044 25172 30100
rect 25340 29932 25396 29988
rect 25116 28642 25172 28644
rect 25116 28590 25118 28642
rect 25118 28590 25170 28642
rect 25170 28590 25172 28642
rect 25116 28588 25172 28590
rect 25900 30380 25956 30436
rect 25564 29596 25620 29652
rect 26236 30994 26292 30996
rect 26236 30942 26238 30994
rect 26238 30942 26290 30994
rect 26290 30942 26292 30994
rect 26236 30940 26292 30942
rect 26012 29986 26068 29988
rect 26012 29934 26014 29986
rect 26014 29934 26066 29986
rect 26066 29934 26068 29986
rect 26012 29932 26068 29934
rect 25676 29260 25732 29316
rect 25340 28082 25396 28084
rect 25340 28030 25342 28082
rect 25342 28030 25394 28082
rect 25394 28030 25396 28082
rect 25340 28028 25396 28030
rect 25228 27858 25284 27860
rect 25228 27806 25230 27858
rect 25230 27806 25282 27858
rect 25282 27806 25284 27858
rect 25228 27804 25284 27806
rect 24220 27132 24276 27188
rect 25452 27580 25508 27636
rect 25452 26236 25508 26292
rect 26012 29148 26068 29204
rect 26012 28642 26068 28644
rect 26012 28590 26014 28642
rect 26014 28590 26066 28642
rect 26066 28590 26068 28642
rect 26012 28588 26068 28590
rect 27356 36876 27412 36932
rect 27132 35586 27188 35588
rect 27132 35534 27134 35586
rect 27134 35534 27186 35586
rect 27186 35534 27188 35586
rect 27132 35532 27188 35534
rect 27132 35308 27188 35364
rect 27020 35084 27076 35140
rect 27132 34972 27188 35028
rect 27580 36594 27636 36596
rect 27580 36542 27582 36594
rect 27582 36542 27634 36594
rect 27634 36542 27636 36594
rect 27580 36540 27636 36542
rect 28364 38162 28420 38164
rect 28364 38110 28366 38162
rect 28366 38110 28418 38162
rect 28418 38110 28420 38162
rect 28364 38108 28420 38110
rect 28700 39900 28756 39956
rect 28588 39116 28644 39172
rect 29148 39900 29204 39956
rect 29820 48242 29876 48244
rect 29820 48190 29822 48242
rect 29822 48190 29874 48242
rect 29874 48190 29876 48242
rect 29820 48188 29876 48190
rect 29596 46844 29652 46900
rect 30716 49980 30772 50036
rect 32396 50370 32452 50372
rect 32396 50318 32398 50370
rect 32398 50318 32450 50370
rect 32450 50318 32452 50370
rect 32396 50316 32452 50318
rect 31836 49644 31892 49700
rect 31724 48524 31780 48580
rect 31500 48354 31556 48356
rect 31500 48302 31502 48354
rect 31502 48302 31554 48354
rect 31554 48302 31556 48354
rect 31500 48300 31556 48302
rect 35196 55690 35252 55692
rect 35196 55638 35198 55690
rect 35198 55638 35250 55690
rect 35250 55638 35252 55690
rect 35196 55636 35252 55638
rect 35300 55690 35356 55692
rect 35300 55638 35302 55690
rect 35302 55638 35354 55690
rect 35354 55638 35356 55690
rect 35300 55636 35356 55638
rect 35404 55690 35460 55692
rect 35404 55638 35406 55690
rect 35406 55638 35458 55690
rect 35458 55638 35460 55690
rect 35404 55636 35460 55638
rect 36316 54572 36372 54628
rect 33964 54348 34020 54404
rect 33628 53788 33684 53844
rect 36316 54402 36372 54404
rect 36316 54350 36318 54402
rect 36318 54350 36370 54402
rect 36370 54350 36372 54402
rect 36316 54348 36372 54350
rect 35196 54122 35252 54124
rect 35196 54070 35198 54122
rect 35198 54070 35250 54122
rect 35250 54070 35252 54122
rect 35196 54068 35252 54070
rect 35300 54122 35356 54124
rect 35300 54070 35302 54122
rect 35302 54070 35354 54122
rect 35354 54070 35356 54122
rect 35300 54068 35356 54070
rect 35404 54122 35460 54124
rect 35404 54070 35406 54122
rect 35406 54070 35458 54122
rect 35458 54070 35460 54122
rect 35404 54068 35460 54070
rect 33964 52946 34020 52948
rect 33964 52894 33966 52946
rect 33966 52894 34018 52946
rect 34018 52894 34020 52946
rect 33964 52892 34020 52894
rect 34412 53116 34468 53172
rect 32956 50316 33012 50372
rect 32172 48300 32228 48356
rect 30940 47964 30996 48020
rect 31500 47852 31556 47908
rect 31276 47458 31332 47460
rect 31276 47406 31278 47458
rect 31278 47406 31330 47458
rect 31330 47406 31332 47458
rect 31276 47404 31332 47406
rect 31164 47180 31220 47236
rect 30380 46508 30436 46564
rect 31164 46620 31220 46676
rect 29596 46396 29652 46452
rect 29372 46060 29428 46116
rect 29372 45276 29428 45332
rect 29372 42754 29428 42756
rect 29372 42702 29374 42754
rect 29374 42702 29426 42754
rect 29426 42702 29428 42754
rect 29372 42700 29428 42702
rect 30156 44492 30212 44548
rect 30044 44268 30100 44324
rect 29932 43372 29988 43428
rect 29596 41970 29652 41972
rect 29596 41918 29598 41970
rect 29598 41918 29650 41970
rect 29650 41918 29652 41970
rect 29596 41916 29652 41918
rect 29596 41186 29652 41188
rect 29596 41134 29598 41186
rect 29598 41134 29650 41186
rect 29650 41134 29652 41186
rect 29596 41132 29652 41134
rect 29372 40124 29428 40180
rect 29484 40572 29540 40628
rect 29484 40236 29540 40292
rect 29260 39564 29316 39620
rect 28588 38220 28644 38276
rect 27916 37154 27972 37156
rect 27916 37102 27918 37154
rect 27918 37102 27970 37154
rect 27970 37102 27972 37154
rect 27916 37100 27972 37102
rect 27916 36876 27972 36932
rect 28028 36316 28084 36372
rect 28028 36092 28084 36148
rect 28588 37100 28644 37156
rect 28700 37884 28756 37940
rect 28476 36428 28532 36484
rect 28364 36370 28420 36372
rect 28364 36318 28366 36370
rect 28366 36318 28418 36370
rect 28418 36318 28420 36370
rect 28364 36316 28420 36318
rect 28476 36258 28532 36260
rect 28476 36206 28478 36258
rect 28478 36206 28530 36258
rect 28530 36206 28532 36258
rect 28476 36204 28532 36206
rect 27020 34076 27076 34132
rect 27020 33292 27076 33348
rect 27020 32620 27076 32676
rect 26796 30156 26852 30212
rect 26684 28812 26740 28868
rect 26348 28754 26404 28756
rect 26348 28702 26350 28754
rect 26350 28702 26402 28754
rect 26402 28702 26404 28754
rect 26348 28700 26404 28702
rect 26684 27858 26740 27860
rect 26684 27806 26686 27858
rect 26686 27806 26738 27858
rect 26738 27806 26740 27858
rect 26684 27804 26740 27806
rect 26460 27692 26516 27748
rect 26908 29148 26964 29204
rect 27244 33628 27300 33684
rect 27356 33292 27412 33348
rect 27580 35420 27636 35476
rect 27804 35698 27860 35700
rect 27804 35646 27806 35698
rect 27806 35646 27858 35698
rect 27858 35646 27860 35698
rect 27804 35644 27860 35646
rect 27804 35308 27860 35364
rect 28028 34690 28084 34692
rect 28028 34638 28030 34690
rect 28030 34638 28082 34690
rect 28082 34638 28084 34690
rect 28028 34636 28084 34638
rect 28476 35420 28532 35476
rect 28252 34300 28308 34356
rect 27580 33906 27636 33908
rect 27580 33854 27582 33906
rect 27582 33854 27634 33906
rect 27634 33854 27636 33906
rect 27580 33852 27636 33854
rect 27804 33628 27860 33684
rect 27692 33122 27748 33124
rect 27692 33070 27694 33122
rect 27694 33070 27746 33122
rect 27746 33070 27748 33122
rect 27692 33068 27748 33070
rect 27580 32732 27636 32788
rect 27132 30882 27188 30884
rect 27132 30830 27134 30882
rect 27134 30830 27186 30882
rect 27186 30830 27188 30882
rect 27132 30828 27188 30830
rect 27132 29650 27188 29652
rect 27132 29598 27134 29650
rect 27134 29598 27186 29650
rect 27186 29598 27188 29650
rect 27132 29596 27188 29598
rect 27692 32562 27748 32564
rect 27692 32510 27694 32562
rect 27694 32510 27746 32562
rect 27746 32510 27748 32562
rect 27692 32508 27748 32510
rect 28028 33346 28084 33348
rect 28028 33294 28030 33346
rect 28030 33294 28082 33346
rect 28082 33294 28084 33346
rect 28028 33292 28084 33294
rect 28028 32732 28084 32788
rect 28252 33234 28308 33236
rect 28252 33182 28254 33234
rect 28254 33182 28306 33234
rect 28306 33182 28308 33234
rect 28252 33180 28308 33182
rect 29708 37826 29764 37828
rect 29708 37774 29710 37826
rect 29710 37774 29762 37826
rect 29762 37774 29764 37826
rect 29708 37772 29764 37774
rect 29372 37660 29428 37716
rect 29036 37378 29092 37380
rect 29036 37326 29038 37378
rect 29038 37326 29090 37378
rect 29090 37326 29092 37378
rect 29036 37324 29092 37326
rect 29036 37100 29092 37156
rect 29596 37490 29652 37492
rect 29596 37438 29598 37490
rect 29598 37438 29650 37490
rect 29650 37438 29652 37490
rect 29596 37436 29652 37438
rect 29484 37378 29540 37380
rect 29484 37326 29486 37378
rect 29486 37326 29538 37378
rect 29538 37326 29540 37378
rect 29484 37324 29540 37326
rect 28812 35698 28868 35700
rect 28812 35646 28814 35698
rect 28814 35646 28866 35698
rect 28866 35646 28868 35698
rect 28812 35644 28868 35646
rect 28588 34972 28644 35028
rect 28700 34690 28756 34692
rect 28700 34638 28702 34690
rect 28702 34638 28754 34690
rect 28754 34638 28756 34690
rect 28700 34636 28756 34638
rect 28812 33292 28868 33348
rect 28364 32674 28420 32676
rect 28364 32622 28366 32674
rect 28366 32622 28418 32674
rect 28418 32622 28420 32674
rect 28364 32620 28420 32622
rect 28924 32508 28980 32564
rect 27804 31218 27860 31220
rect 27804 31166 27806 31218
rect 27806 31166 27858 31218
rect 27858 31166 27860 31218
rect 27804 31164 27860 31166
rect 27692 30492 27748 30548
rect 28028 30828 28084 30884
rect 28028 30268 28084 30324
rect 28364 30380 28420 30436
rect 27580 30156 27636 30212
rect 27244 28812 27300 28868
rect 27356 29260 27412 29316
rect 27356 28754 27412 28756
rect 27356 28702 27358 28754
rect 27358 28702 27410 28754
rect 27410 28702 27412 28754
rect 27356 28700 27412 28702
rect 27356 27970 27412 27972
rect 27356 27918 27358 27970
rect 27358 27918 27410 27970
rect 27410 27918 27412 27970
rect 27356 27916 27412 27918
rect 26796 26236 26852 26292
rect 27916 29932 27972 29988
rect 27692 29650 27748 29652
rect 27692 29598 27694 29650
rect 27694 29598 27746 29650
rect 27746 29598 27748 29650
rect 27692 29596 27748 29598
rect 27804 29314 27860 29316
rect 27804 29262 27806 29314
rect 27806 29262 27858 29314
rect 27858 29262 27860 29314
rect 27804 29260 27860 29262
rect 28364 29426 28420 29428
rect 28364 29374 28366 29426
rect 28366 29374 28418 29426
rect 28418 29374 28420 29426
rect 28364 29372 28420 29374
rect 25564 26124 25620 26180
rect 24444 25788 24500 25844
rect 25340 25564 25396 25620
rect 24444 25116 24500 25172
rect 24220 24668 24276 24724
rect 25788 24946 25844 24948
rect 25788 24894 25790 24946
rect 25790 24894 25842 24946
rect 25842 24894 25844 24946
rect 25788 24892 25844 24894
rect 24108 24556 24164 24612
rect 24332 24220 24388 24276
rect 25004 24668 25060 24724
rect 24444 23996 24500 24052
rect 25228 24610 25284 24612
rect 25228 24558 25230 24610
rect 25230 24558 25282 24610
rect 25282 24558 25284 24610
rect 25228 24556 25284 24558
rect 24780 23938 24836 23940
rect 24780 23886 24782 23938
rect 24782 23886 24834 23938
rect 24834 23886 24836 23938
rect 24780 23884 24836 23886
rect 26236 24946 26292 24948
rect 26236 24894 26238 24946
rect 26238 24894 26290 24946
rect 26290 24894 26292 24946
rect 26236 24892 26292 24894
rect 25788 24050 25844 24052
rect 25788 23998 25790 24050
rect 25790 23998 25842 24050
rect 25842 23998 25844 24050
rect 25788 23996 25844 23998
rect 25452 23884 25508 23940
rect 23996 23436 24052 23492
rect 22204 23378 22260 23380
rect 22204 23326 22206 23378
rect 22206 23326 22258 23378
rect 22258 23326 22260 23378
rect 22204 23324 22260 23326
rect 22988 23378 23044 23380
rect 22988 23326 22990 23378
rect 22990 23326 23042 23378
rect 23042 23326 23044 23378
rect 22988 23324 23044 23326
rect 21308 23266 21364 23268
rect 21308 23214 21310 23266
rect 21310 23214 21362 23266
rect 21362 23214 21364 23266
rect 21308 23212 21364 23214
rect 28252 28700 28308 28756
rect 27804 26572 27860 26628
rect 28476 28700 28532 28756
rect 27916 27804 27972 27860
rect 27132 25618 27188 25620
rect 27132 25566 27134 25618
rect 27134 25566 27186 25618
rect 27186 25566 27188 25618
rect 27132 25564 27188 25566
rect 27020 23100 27076 23156
rect 27804 25282 27860 25284
rect 27804 25230 27806 25282
rect 27806 25230 27858 25282
rect 27858 25230 27860 25282
rect 27804 25228 27860 25230
rect 28140 27746 28196 27748
rect 28140 27694 28142 27746
rect 28142 27694 28194 27746
rect 28194 27694 28196 27746
rect 28140 27692 28196 27694
rect 28700 30380 28756 30436
rect 28924 29372 28980 29428
rect 29260 36258 29316 36260
rect 29260 36206 29262 36258
rect 29262 36206 29314 36258
rect 29314 36206 29316 36258
rect 29260 36204 29316 36206
rect 29260 35084 29316 35140
rect 29372 35196 29428 35252
rect 29260 34354 29316 34356
rect 29260 34302 29262 34354
rect 29262 34302 29314 34354
rect 29314 34302 29316 34354
rect 29260 34300 29316 34302
rect 29260 33234 29316 33236
rect 29260 33182 29262 33234
rect 29262 33182 29314 33234
rect 29314 33182 29316 33234
rect 29260 33180 29316 33182
rect 29148 33068 29204 33124
rect 30828 44322 30884 44324
rect 30828 44270 30830 44322
rect 30830 44270 30882 44322
rect 30882 44270 30884 44322
rect 30828 44268 30884 44270
rect 30604 43708 30660 43764
rect 31052 43372 31108 43428
rect 30268 42476 30324 42532
rect 30828 42140 30884 42196
rect 30156 41916 30212 41972
rect 31052 41074 31108 41076
rect 31052 41022 31054 41074
rect 31054 41022 31106 41074
rect 31106 41022 31108 41074
rect 31052 41020 31108 41022
rect 30380 40962 30436 40964
rect 30380 40910 30382 40962
rect 30382 40910 30434 40962
rect 30434 40910 30436 40962
rect 30380 40908 30436 40910
rect 30044 40796 30100 40852
rect 30156 40402 30212 40404
rect 30156 40350 30158 40402
rect 30158 40350 30210 40402
rect 30210 40350 30212 40402
rect 30156 40348 30212 40350
rect 30828 40236 30884 40292
rect 32060 47570 32116 47572
rect 32060 47518 32062 47570
rect 32062 47518 32114 47570
rect 32114 47518 32116 47570
rect 32060 47516 32116 47518
rect 31948 47292 32004 47348
rect 31836 45890 31892 45892
rect 31836 45838 31838 45890
rect 31838 45838 31890 45890
rect 31890 45838 31892 45890
rect 31836 45836 31892 45838
rect 31724 44156 31780 44212
rect 31724 43650 31780 43652
rect 31724 43598 31726 43650
rect 31726 43598 31778 43650
rect 31778 43598 31780 43650
rect 31724 43596 31780 43598
rect 32060 46002 32116 46004
rect 32060 45950 32062 46002
rect 32062 45950 32114 46002
rect 32114 45950 32116 46002
rect 32060 45948 32116 45950
rect 34524 53564 34580 53620
rect 37100 55020 37156 55076
rect 36988 53676 37044 53732
rect 36764 53058 36820 53060
rect 36764 53006 36766 53058
rect 36766 53006 36818 53058
rect 36818 53006 36820 53058
rect 36764 53004 36820 53006
rect 36540 52780 36596 52836
rect 35196 52554 35252 52556
rect 35196 52502 35198 52554
rect 35198 52502 35250 52554
rect 35250 52502 35252 52554
rect 35196 52500 35252 52502
rect 35300 52554 35356 52556
rect 35300 52502 35302 52554
rect 35302 52502 35354 52554
rect 35354 52502 35356 52554
rect 35300 52500 35356 52502
rect 35404 52554 35460 52556
rect 35404 52502 35406 52554
rect 35406 52502 35458 52554
rect 35458 52502 35460 52554
rect 35404 52500 35460 52502
rect 35196 50986 35252 50988
rect 35196 50934 35198 50986
rect 35198 50934 35250 50986
rect 35250 50934 35252 50986
rect 35196 50932 35252 50934
rect 35300 50986 35356 50988
rect 35300 50934 35302 50986
rect 35302 50934 35354 50986
rect 35354 50934 35356 50986
rect 35300 50932 35356 50934
rect 35404 50986 35460 50988
rect 35404 50934 35406 50986
rect 35406 50934 35458 50986
rect 35458 50934 35460 50986
rect 35404 50932 35460 50934
rect 37100 50652 37156 50708
rect 33516 50316 33572 50372
rect 33068 50034 33124 50036
rect 33068 49982 33070 50034
rect 33070 49982 33122 50034
rect 33122 49982 33124 50034
rect 33068 49980 33124 49982
rect 34076 49980 34132 50036
rect 33292 49810 33348 49812
rect 33292 49758 33294 49810
rect 33294 49758 33346 49810
rect 33346 49758 33348 49810
rect 33292 49756 33348 49758
rect 33180 49698 33236 49700
rect 33180 49646 33182 49698
rect 33182 49646 33234 49698
rect 33234 49646 33236 49698
rect 33180 49644 33236 49646
rect 33516 48636 33572 48692
rect 33068 48524 33124 48580
rect 32844 48076 32900 48132
rect 32844 47404 32900 47460
rect 33180 47458 33236 47460
rect 33180 47406 33182 47458
rect 33182 47406 33234 47458
rect 33234 47406 33236 47458
rect 33180 47404 33236 47406
rect 33292 47068 33348 47124
rect 33964 49532 34020 49588
rect 32620 46674 32676 46676
rect 32620 46622 32622 46674
rect 32622 46622 32674 46674
rect 32674 46622 32676 46674
rect 32620 46620 32676 46622
rect 32732 46844 32788 46900
rect 32508 46508 32564 46564
rect 33292 46674 33348 46676
rect 33292 46622 33294 46674
rect 33294 46622 33346 46674
rect 33346 46622 33348 46674
rect 33292 46620 33348 46622
rect 32956 46396 33012 46452
rect 33628 47180 33684 47236
rect 33740 46956 33796 47012
rect 33516 45724 33572 45780
rect 34300 49532 34356 49588
rect 34188 48636 34244 48692
rect 34076 46844 34132 46900
rect 37100 50316 37156 50372
rect 34860 49698 34916 49700
rect 34860 49646 34862 49698
rect 34862 49646 34914 49698
rect 34914 49646 34916 49698
rect 34860 49644 34916 49646
rect 34748 49532 34804 49588
rect 34972 47458 35028 47460
rect 34972 47406 34974 47458
rect 34974 47406 35026 47458
rect 35026 47406 35028 47458
rect 34972 47404 35028 47406
rect 35420 49532 35476 49588
rect 35644 49644 35700 49700
rect 35196 49418 35252 49420
rect 35196 49366 35198 49418
rect 35198 49366 35250 49418
rect 35250 49366 35252 49418
rect 35196 49364 35252 49366
rect 35300 49418 35356 49420
rect 35300 49366 35302 49418
rect 35302 49366 35354 49418
rect 35354 49366 35356 49418
rect 35300 49364 35356 49366
rect 35404 49418 35460 49420
rect 35404 49366 35406 49418
rect 35406 49366 35458 49418
rect 35458 49366 35460 49418
rect 35404 49364 35460 49366
rect 36428 48748 36484 48804
rect 37100 48636 37156 48692
rect 37772 55074 37828 55076
rect 37772 55022 37774 55074
rect 37774 55022 37826 55074
rect 37826 55022 37828 55074
rect 37772 55020 37828 55022
rect 38892 55804 38948 55860
rect 43260 56252 43316 56308
rect 44604 56306 44660 56308
rect 44604 56254 44606 56306
rect 44606 56254 44658 56306
rect 44658 56254 44660 56306
rect 44604 56252 44660 56254
rect 40460 55804 40516 55860
rect 38220 54572 38276 54628
rect 39900 55074 39956 55076
rect 39900 55022 39902 55074
rect 39902 55022 39954 55074
rect 39954 55022 39956 55074
rect 39900 55020 39956 55022
rect 40348 55020 40404 55076
rect 39116 54684 39172 54740
rect 40348 54738 40404 54740
rect 40348 54686 40350 54738
rect 40350 54686 40402 54738
rect 40402 54686 40404 54738
rect 40348 54684 40404 54686
rect 40796 54684 40852 54740
rect 38892 54626 38948 54628
rect 38892 54574 38894 54626
rect 38894 54574 38946 54626
rect 38946 54574 38948 54626
rect 38892 54572 38948 54574
rect 37884 54236 37940 54292
rect 39452 53900 39508 53956
rect 39116 53788 39172 53844
rect 38444 53564 38500 53620
rect 37772 52946 37828 52948
rect 37772 52894 37774 52946
rect 37774 52894 37826 52946
rect 37826 52894 37828 52946
rect 37772 52892 37828 52894
rect 37660 52834 37716 52836
rect 37660 52782 37662 52834
rect 37662 52782 37714 52834
rect 37714 52782 37716 52834
rect 37660 52780 37716 52782
rect 37436 52108 37492 52164
rect 38332 52162 38388 52164
rect 38332 52110 38334 52162
rect 38334 52110 38386 52162
rect 38386 52110 38388 52162
rect 38332 52108 38388 52110
rect 38108 51660 38164 51716
rect 39228 52050 39284 52052
rect 39228 51998 39230 52050
rect 39230 51998 39282 52050
rect 39282 51998 39284 52050
rect 39228 51996 39284 51998
rect 38668 51548 38724 51604
rect 37324 51436 37380 51492
rect 35196 47850 35252 47852
rect 35196 47798 35198 47850
rect 35198 47798 35250 47850
rect 35250 47798 35252 47850
rect 35196 47796 35252 47798
rect 35300 47850 35356 47852
rect 35300 47798 35302 47850
rect 35302 47798 35354 47850
rect 35354 47798 35356 47850
rect 35300 47796 35356 47798
rect 35404 47850 35460 47852
rect 35404 47798 35406 47850
rect 35406 47798 35458 47850
rect 35458 47798 35460 47850
rect 35404 47796 35460 47798
rect 35756 47740 35812 47796
rect 38444 51378 38500 51380
rect 38444 51326 38446 51378
rect 38446 51326 38498 51378
rect 38498 51326 38500 51378
rect 38444 51324 38500 51326
rect 37884 51212 37940 51268
rect 38780 51378 38836 51380
rect 38780 51326 38782 51378
rect 38782 51326 38834 51378
rect 38834 51326 38836 51378
rect 38780 51324 38836 51326
rect 38892 51266 38948 51268
rect 38892 51214 38894 51266
rect 38894 51214 38946 51266
rect 38946 51214 38948 51266
rect 38892 51212 38948 51214
rect 38444 51100 38500 51156
rect 39004 51100 39060 51156
rect 39228 51154 39284 51156
rect 39228 51102 39230 51154
rect 39230 51102 39282 51154
rect 39282 51102 39284 51154
rect 39228 51100 39284 51102
rect 38556 48636 38612 48692
rect 37324 47740 37380 47796
rect 38332 47740 38388 47796
rect 33404 45612 33460 45668
rect 32172 44492 32228 44548
rect 32732 44380 32788 44436
rect 32956 44210 33012 44212
rect 32956 44158 32958 44210
rect 32958 44158 33010 44210
rect 33010 44158 33012 44210
rect 32956 44156 33012 44158
rect 32620 43650 32676 43652
rect 32620 43598 32622 43650
rect 32622 43598 32674 43650
rect 32674 43598 32676 43650
rect 32620 43596 32676 43598
rect 33292 44156 33348 44212
rect 33516 44268 33572 44324
rect 33068 43650 33124 43652
rect 33068 43598 33070 43650
rect 33070 43598 33122 43650
rect 33122 43598 33124 43650
rect 33068 43596 33124 43598
rect 33404 43650 33460 43652
rect 33404 43598 33406 43650
rect 33406 43598 33458 43650
rect 33458 43598 33460 43650
rect 33404 43596 33460 43598
rect 33516 43260 33572 43316
rect 33516 42754 33572 42756
rect 33516 42702 33518 42754
rect 33518 42702 33570 42754
rect 33570 42702 33572 42754
rect 33516 42700 33572 42702
rect 32844 42530 32900 42532
rect 32844 42478 32846 42530
rect 32846 42478 32898 42530
rect 32898 42478 32900 42530
rect 32844 42476 32900 42478
rect 32060 41916 32116 41972
rect 32844 42028 32900 42084
rect 33964 42364 34020 42420
rect 33516 41970 33572 41972
rect 33516 41918 33518 41970
rect 33518 41918 33570 41970
rect 33570 41918 33572 41970
rect 33516 41916 33572 41918
rect 34188 45724 34244 45780
rect 34524 46172 34580 46228
rect 37772 47628 37828 47684
rect 35756 47404 35812 47460
rect 38108 47458 38164 47460
rect 38108 47406 38110 47458
rect 38110 47406 38162 47458
rect 38162 47406 38164 47458
rect 38108 47404 38164 47406
rect 35084 47180 35140 47236
rect 34860 46844 34916 46900
rect 35196 46732 35252 46788
rect 36652 46786 36708 46788
rect 36652 46734 36654 46786
rect 36654 46734 36706 46786
rect 36706 46734 36708 46786
rect 36652 46732 36708 46734
rect 35196 46282 35252 46284
rect 35196 46230 35198 46282
rect 35198 46230 35250 46282
rect 35250 46230 35252 46282
rect 35196 46228 35252 46230
rect 35300 46282 35356 46284
rect 35300 46230 35302 46282
rect 35302 46230 35354 46282
rect 35354 46230 35356 46282
rect 35300 46228 35356 46230
rect 35404 46282 35460 46284
rect 35404 46230 35406 46282
rect 35406 46230 35458 46282
rect 35458 46230 35460 46282
rect 35404 46228 35460 46230
rect 34188 44322 34244 44324
rect 34188 44270 34190 44322
rect 34190 44270 34242 44322
rect 34242 44270 34244 44322
rect 34188 44268 34244 44270
rect 34412 42924 34468 42980
rect 34524 45612 34580 45668
rect 37548 44940 37604 44996
rect 35196 44714 35252 44716
rect 35196 44662 35198 44714
rect 35198 44662 35250 44714
rect 35250 44662 35252 44714
rect 35196 44660 35252 44662
rect 35300 44714 35356 44716
rect 35300 44662 35302 44714
rect 35302 44662 35354 44714
rect 35354 44662 35356 44714
rect 35300 44660 35356 44662
rect 35404 44714 35460 44716
rect 35404 44662 35406 44714
rect 35406 44662 35458 44714
rect 35458 44662 35460 44714
rect 35404 44660 35460 44662
rect 34748 44492 34804 44548
rect 35420 44492 35476 44548
rect 36316 44268 36372 44324
rect 34972 43596 35028 43652
rect 34076 41858 34132 41860
rect 34076 41806 34078 41858
rect 34078 41806 34130 41858
rect 34130 41806 34132 41858
rect 34076 41804 34132 41806
rect 35196 43146 35252 43148
rect 35196 43094 35198 43146
rect 35198 43094 35250 43146
rect 35250 43094 35252 43146
rect 35196 43092 35252 43094
rect 35300 43146 35356 43148
rect 35300 43094 35302 43146
rect 35302 43094 35354 43146
rect 35354 43094 35356 43146
rect 35300 43092 35356 43094
rect 35404 43146 35460 43148
rect 35404 43094 35406 43146
rect 35406 43094 35458 43146
rect 35458 43094 35460 43146
rect 35404 43092 35460 43094
rect 35308 42924 35364 42980
rect 34636 42028 34692 42084
rect 34524 41916 34580 41972
rect 33516 41186 33572 41188
rect 33516 41134 33518 41186
rect 33518 41134 33570 41186
rect 33570 41134 33572 41186
rect 33516 41132 33572 41134
rect 31276 40460 31332 40516
rect 30044 39618 30100 39620
rect 30044 39566 30046 39618
rect 30046 39566 30098 39618
rect 30098 39566 30100 39618
rect 30044 39564 30100 39566
rect 30044 38162 30100 38164
rect 30044 38110 30046 38162
rect 30046 38110 30098 38162
rect 30098 38110 30100 38162
rect 30044 38108 30100 38110
rect 30044 37100 30100 37156
rect 29932 36764 29988 36820
rect 29708 36258 29764 36260
rect 29708 36206 29710 36258
rect 29710 36206 29762 36258
rect 29762 36206 29764 36258
rect 29708 36204 29764 36206
rect 29820 35196 29876 35252
rect 29708 34972 29764 35028
rect 30268 39842 30324 39844
rect 30268 39790 30270 39842
rect 30270 39790 30322 39842
rect 30322 39790 30324 39842
rect 30268 39788 30324 39790
rect 31052 39340 31108 39396
rect 30492 38050 30548 38052
rect 30492 37998 30494 38050
rect 30494 37998 30546 38050
rect 30546 37998 30548 38050
rect 30492 37996 30548 37998
rect 30604 37938 30660 37940
rect 30604 37886 30606 37938
rect 30606 37886 30658 37938
rect 30658 37886 30660 37938
rect 30604 37884 30660 37886
rect 30492 37042 30548 37044
rect 30492 36990 30494 37042
rect 30494 36990 30546 37042
rect 30546 36990 30548 37042
rect 30492 36988 30548 36990
rect 30380 34636 30436 34692
rect 30268 34018 30324 34020
rect 30268 33966 30270 34018
rect 30270 33966 30322 34018
rect 30322 33966 30324 34018
rect 30268 33964 30324 33966
rect 29484 32508 29540 32564
rect 29372 31164 29428 31220
rect 29708 31554 29764 31556
rect 29708 31502 29710 31554
rect 29710 31502 29762 31554
rect 29762 31502 29764 31554
rect 29708 31500 29764 31502
rect 29708 31164 29764 31220
rect 29260 29986 29316 29988
rect 29260 29934 29262 29986
rect 29262 29934 29314 29986
rect 29314 29934 29316 29986
rect 29260 29932 29316 29934
rect 29148 28700 29204 28756
rect 29596 29260 29652 29316
rect 28700 28364 28756 28420
rect 29708 29372 29764 29428
rect 30716 34636 30772 34692
rect 30268 29596 30324 29652
rect 30492 30044 30548 30100
rect 30492 29148 30548 29204
rect 29260 28364 29316 28420
rect 29708 28082 29764 28084
rect 29708 28030 29710 28082
rect 29710 28030 29762 28082
rect 29762 28030 29764 28082
rect 29708 28028 29764 28030
rect 30604 28082 30660 28084
rect 30604 28030 30606 28082
rect 30606 28030 30658 28082
rect 30658 28030 30660 28082
rect 30604 28028 30660 28030
rect 30044 27858 30100 27860
rect 30044 27806 30046 27858
rect 30046 27806 30098 27858
rect 30098 27806 30100 27858
rect 30044 27804 30100 27806
rect 28588 27244 28644 27300
rect 29148 27244 29204 27300
rect 32172 40348 32228 40404
rect 31388 39228 31444 39284
rect 31164 38444 31220 38500
rect 31276 38108 31332 38164
rect 31052 37996 31108 38052
rect 30940 35980 30996 36036
rect 30940 35196 30996 35252
rect 30940 31554 30996 31556
rect 30940 31502 30942 31554
rect 30942 31502 30994 31554
rect 30994 31502 30996 31554
rect 30940 31500 30996 31502
rect 30940 30210 30996 30212
rect 30940 30158 30942 30210
rect 30942 30158 30994 30210
rect 30994 30158 30996 30210
rect 30940 30156 30996 30158
rect 31500 37436 31556 37492
rect 32844 39452 32900 39508
rect 32060 37938 32116 37940
rect 32060 37886 32062 37938
rect 32062 37886 32114 37938
rect 32114 37886 32116 37938
rect 32060 37884 32116 37886
rect 31724 37772 31780 37828
rect 32172 37772 32228 37828
rect 31724 37436 31780 37492
rect 32060 37490 32116 37492
rect 32060 37438 32062 37490
rect 32062 37438 32114 37490
rect 32114 37438 32116 37490
rect 32060 37436 32116 37438
rect 32396 38444 32452 38500
rect 32844 37996 32900 38052
rect 32396 37212 32452 37268
rect 32732 37772 32788 37828
rect 31948 37154 32004 37156
rect 31948 37102 31950 37154
rect 31950 37102 32002 37154
rect 32002 37102 32004 37154
rect 31948 37100 32004 37102
rect 31612 35084 31668 35140
rect 31724 35644 31780 35700
rect 32284 35644 32340 35700
rect 31724 34748 31780 34804
rect 31388 33516 31444 33572
rect 32172 33570 32228 33572
rect 32172 33518 32174 33570
rect 32174 33518 32226 33570
rect 32226 33518 32228 33570
rect 32172 33516 32228 33518
rect 32396 33516 32452 33572
rect 32172 32732 32228 32788
rect 31500 30322 31556 30324
rect 31500 30270 31502 30322
rect 31502 30270 31554 30322
rect 31554 30270 31556 30322
rect 31500 30268 31556 30270
rect 31948 30210 32004 30212
rect 31948 30158 31950 30210
rect 31950 30158 32002 30210
rect 32002 30158 32004 30210
rect 31948 30156 32004 30158
rect 31052 30044 31108 30100
rect 30828 28140 30884 28196
rect 33068 40962 33124 40964
rect 33068 40910 33070 40962
rect 33070 40910 33122 40962
rect 33122 40910 33124 40962
rect 33068 40908 33124 40910
rect 34076 40684 34132 40740
rect 34636 41746 34692 41748
rect 34636 41694 34638 41746
rect 34638 41694 34690 41746
rect 34690 41694 34692 41746
rect 34636 41692 34692 41694
rect 35196 42082 35252 42084
rect 35196 42030 35198 42082
rect 35198 42030 35250 42082
rect 35250 42030 35252 42082
rect 35196 42028 35252 42030
rect 35084 41804 35140 41860
rect 34524 40684 34580 40740
rect 34636 40572 34692 40628
rect 35420 41916 35476 41972
rect 35196 41578 35252 41580
rect 35196 41526 35198 41578
rect 35198 41526 35250 41578
rect 35250 41526 35252 41578
rect 35196 41524 35252 41526
rect 35300 41578 35356 41580
rect 35300 41526 35302 41578
rect 35302 41526 35354 41578
rect 35354 41526 35356 41578
rect 35300 41524 35356 41526
rect 35404 41578 35460 41580
rect 35404 41526 35406 41578
rect 35406 41526 35458 41578
rect 35458 41526 35460 41578
rect 35404 41524 35460 41526
rect 35308 41410 35364 41412
rect 35308 41358 35310 41410
rect 35310 41358 35362 41410
rect 35362 41358 35364 41410
rect 35308 41356 35364 41358
rect 35308 40572 35364 40628
rect 35308 40402 35364 40404
rect 35308 40350 35310 40402
rect 35310 40350 35362 40402
rect 35362 40350 35364 40402
rect 35308 40348 35364 40350
rect 35644 41356 35700 41412
rect 35756 41692 35812 41748
rect 35196 40236 35252 40292
rect 35532 40124 35588 40180
rect 35196 40010 35252 40012
rect 35196 39958 35198 40010
rect 35198 39958 35250 40010
rect 35250 39958 35252 40010
rect 35196 39956 35252 39958
rect 35300 40010 35356 40012
rect 35300 39958 35302 40010
rect 35302 39958 35354 40010
rect 35354 39958 35356 40010
rect 35300 39956 35356 39958
rect 35404 40010 35460 40012
rect 35404 39958 35406 40010
rect 35406 39958 35458 40010
rect 35458 39958 35460 40010
rect 35404 39956 35460 39958
rect 33740 39506 33796 39508
rect 33740 39454 33742 39506
rect 33742 39454 33794 39506
rect 33794 39454 33796 39506
rect 33740 39452 33796 39454
rect 33628 39228 33684 39284
rect 34300 38668 34356 38724
rect 34188 38162 34244 38164
rect 34188 38110 34190 38162
rect 34190 38110 34242 38162
rect 34242 38110 34244 38162
rect 34188 38108 34244 38110
rect 33292 37884 33348 37940
rect 33180 36482 33236 36484
rect 33180 36430 33182 36482
rect 33182 36430 33234 36482
rect 33234 36430 33236 36482
rect 33180 36428 33236 36430
rect 33180 35084 33236 35140
rect 32620 31612 32676 31668
rect 33740 37826 33796 37828
rect 33740 37774 33742 37826
rect 33742 37774 33794 37826
rect 33794 37774 33796 37826
rect 33740 37772 33796 37774
rect 34188 37266 34244 37268
rect 34188 37214 34190 37266
rect 34190 37214 34242 37266
rect 34242 37214 34244 37266
rect 34188 37212 34244 37214
rect 33852 36258 33908 36260
rect 33852 36206 33854 36258
rect 33854 36206 33906 36258
rect 33906 36206 33908 36258
rect 33852 36204 33908 36206
rect 34412 35868 34468 35924
rect 33404 35196 33460 35252
rect 34636 38668 34692 38724
rect 33292 33516 33348 33572
rect 33180 33404 33236 33460
rect 33852 33234 33908 33236
rect 33852 33182 33854 33234
rect 33854 33182 33906 33234
rect 33906 33182 33908 33234
rect 33852 33180 33908 33182
rect 33404 32620 33460 32676
rect 33852 32956 33908 33012
rect 33180 31218 33236 31220
rect 33180 31166 33182 31218
rect 33182 31166 33234 31218
rect 33234 31166 33236 31218
rect 33180 31164 33236 31166
rect 33740 30940 33796 30996
rect 32844 29932 32900 29988
rect 34188 32508 34244 32564
rect 34300 33516 34356 33572
rect 34188 31052 34244 31108
rect 35084 38668 35140 38724
rect 35196 38442 35252 38444
rect 35196 38390 35198 38442
rect 35198 38390 35250 38442
rect 35250 38390 35252 38442
rect 35196 38388 35252 38390
rect 35300 38442 35356 38444
rect 35300 38390 35302 38442
rect 35302 38390 35354 38442
rect 35354 38390 35356 38442
rect 35300 38388 35356 38390
rect 35404 38442 35460 38444
rect 35404 38390 35406 38442
rect 35406 38390 35458 38442
rect 35458 38390 35460 38442
rect 35404 38388 35460 38390
rect 35196 36874 35252 36876
rect 35196 36822 35198 36874
rect 35198 36822 35250 36874
rect 35250 36822 35252 36874
rect 35196 36820 35252 36822
rect 35300 36874 35356 36876
rect 35300 36822 35302 36874
rect 35302 36822 35354 36874
rect 35354 36822 35356 36874
rect 35300 36820 35356 36822
rect 35404 36874 35460 36876
rect 35404 36822 35406 36874
rect 35406 36822 35458 36874
rect 35458 36822 35460 36874
rect 35404 36820 35460 36822
rect 36092 40684 36148 40740
rect 40012 51602 40068 51604
rect 40012 51550 40014 51602
rect 40014 51550 40066 51602
rect 40066 51550 40068 51602
rect 40012 51548 40068 51550
rect 40348 50988 40404 51044
rect 40012 48636 40068 48692
rect 39452 48188 39508 48244
rect 38780 47180 38836 47236
rect 38892 47404 38948 47460
rect 38444 46732 38500 46788
rect 38668 46956 38724 47012
rect 38556 45890 38612 45892
rect 38556 45838 38558 45890
rect 38558 45838 38610 45890
rect 38610 45838 38612 45890
rect 38556 45836 38612 45838
rect 39228 46956 39284 47012
rect 39116 46844 39172 46900
rect 39452 45052 39508 45108
rect 39564 46732 39620 46788
rect 38556 44268 38612 44324
rect 37436 44210 37492 44212
rect 37436 44158 37438 44210
rect 37438 44158 37490 44210
rect 37490 44158 37492 44210
rect 37436 44156 37492 44158
rect 36988 43484 37044 43540
rect 36316 40348 36372 40404
rect 36428 43260 36484 43316
rect 35756 38892 35812 38948
rect 35868 40236 35924 40292
rect 36428 40124 36484 40180
rect 37212 43426 37268 43428
rect 37212 43374 37214 43426
rect 37214 43374 37266 43426
rect 37266 43374 37268 43426
rect 37212 43372 37268 43374
rect 38668 43372 38724 43428
rect 38668 42866 38724 42868
rect 38668 42814 38670 42866
rect 38670 42814 38722 42866
rect 38722 42814 38724 42866
rect 38668 42812 38724 42814
rect 39116 44322 39172 44324
rect 39116 44270 39118 44322
rect 39118 44270 39170 44322
rect 39170 44270 39172 44322
rect 39116 44268 39172 44270
rect 39452 43596 39508 43652
rect 39228 42812 39284 42868
rect 38556 42754 38612 42756
rect 38556 42702 38558 42754
rect 38558 42702 38610 42754
rect 38610 42702 38612 42754
rect 38556 42700 38612 42702
rect 39004 42642 39060 42644
rect 39004 42590 39006 42642
rect 39006 42590 39058 42642
rect 39058 42590 39060 42642
rect 39004 42588 39060 42590
rect 39788 46956 39844 47012
rect 40012 47404 40068 47460
rect 40460 50706 40516 50708
rect 40460 50654 40462 50706
rect 40462 50654 40514 50706
rect 40514 50654 40516 50706
rect 40460 50652 40516 50654
rect 40348 46956 40404 47012
rect 41356 54684 41412 54740
rect 41244 54572 41300 54628
rect 40908 54460 40964 54516
rect 41020 53170 41076 53172
rect 41020 53118 41022 53170
rect 41022 53118 41074 53170
rect 41074 53118 41076 53170
rect 41020 53116 41076 53118
rect 41692 54626 41748 54628
rect 41692 54574 41694 54626
rect 41694 54574 41746 54626
rect 41746 54574 41748 54626
rect 41692 54572 41748 54574
rect 41692 53788 41748 53844
rect 41244 53730 41300 53732
rect 41244 53678 41246 53730
rect 41246 53678 41298 53730
rect 41298 53678 41300 53730
rect 41244 53676 41300 53678
rect 41580 53004 41636 53060
rect 41468 52892 41524 52948
rect 41916 53004 41972 53060
rect 47740 56252 47796 56308
rect 48972 56306 49028 56308
rect 48972 56254 48974 56306
rect 48974 56254 49026 56306
rect 49026 56254 49028 56306
rect 48972 56252 49028 56254
rect 50556 56474 50612 56476
rect 50556 56422 50558 56474
rect 50558 56422 50610 56474
rect 50610 56422 50612 56474
rect 50556 56420 50612 56422
rect 50660 56474 50716 56476
rect 50660 56422 50662 56474
rect 50662 56422 50714 56474
rect 50714 56422 50716 56474
rect 50660 56420 50716 56422
rect 50764 56474 50820 56476
rect 50764 56422 50766 56474
rect 50766 56422 50818 56474
rect 50818 56422 50820 56474
rect 50764 56420 50820 56422
rect 49980 56252 50036 56308
rect 52220 56306 52276 56308
rect 52220 56254 52222 56306
rect 52222 56254 52274 56306
rect 52274 56254 52276 56306
rect 52220 56252 52276 56254
rect 45500 55356 45556 55412
rect 46732 55410 46788 55412
rect 46732 55358 46734 55410
rect 46734 55358 46786 55410
rect 46786 55358 46788 55410
rect 46732 55356 46788 55358
rect 43484 53900 43540 53956
rect 43148 53676 43204 53732
rect 41020 51324 41076 51380
rect 41244 51490 41300 51492
rect 41244 51438 41246 51490
rect 41246 51438 41298 51490
rect 41298 51438 41300 51490
rect 41244 51436 41300 51438
rect 40908 50706 40964 50708
rect 40908 50654 40910 50706
rect 40910 50654 40962 50706
rect 40962 50654 40964 50706
rect 40908 50652 40964 50654
rect 42252 52050 42308 52052
rect 42252 51998 42254 52050
rect 42254 51998 42306 52050
rect 42306 51998 42308 52050
rect 42252 51996 42308 51998
rect 41580 51154 41636 51156
rect 41580 51102 41582 51154
rect 41582 51102 41634 51154
rect 41634 51102 41636 51154
rect 41580 51100 41636 51102
rect 42700 52946 42756 52948
rect 42700 52894 42702 52946
rect 42702 52894 42754 52946
rect 42754 52894 42756 52946
rect 42700 52892 42756 52894
rect 42588 52780 42644 52836
rect 42252 51602 42308 51604
rect 42252 51550 42254 51602
rect 42254 51550 42306 51602
rect 42306 51550 42308 51602
rect 42252 51548 42308 51550
rect 44604 53788 44660 53844
rect 41244 50652 41300 50708
rect 42476 50652 42532 50708
rect 44156 50706 44212 50708
rect 44156 50654 44158 50706
rect 44158 50654 44210 50706
rect 44210 50654 44212 50706
rect 44156 50652 44212 50654
rect 42700 47458 42756 47460
rect 42700 47406 42702 47458
rect 42702 47406 42754 47458
rect 42754 47406 42756 47458
rect 42700 47404 42756 47406
rect 41244 47292 41300 47348
rect 41132 46956 41188 47012
rect 40908 46844 40964 46900
rect 42028 47346 42084 47348
rect 42028 47294 42030 47346
rect 42030 47294 42082 47346
rect 42082 47294 42084 47346
rect 42028 47292 42084 47294
rect 41468 46786 41524 46788
rect 41468 46734 41470 46786
rect 41470 46734 41522 46786
rect 41522 46734 41524 46786
rect 41468 46732 41524 46734
rect 40236 45724 40292 45780
rect 40124 44940 40180 44996
rect 40348 45106 40404 45108
rect 40348 45054 40350 45106
rect 40350 45054 40402 45106
rect 40402 45054 40404 45106
rect 40348 45052 40404 45054
rect 41356 45778 41412 45780
rect 41356 45726 41358 45778
rect 41358 45726 41410 45778
rect 41410 45726 41412 45778
rect 41356 45724 41412 45726
rect 40796 44492 40852 44548
rect 39676 43596 39732 43652
rect 40012 43538 40068 43540
rect 40012 43486 40014 43538
rect 40014 43486 40066 43538
rect 40066 43486 40068 43538
rect 40012 43484 40068 43486
rect 40236 43372 40292 43428
rect 41020 43484 41076 43540
rect 41132 43372 41188 43428
rect 44492 44994 44548 44996
rect 44492 44942 44494 44994
rect 44494 44942 44546 44994
rect 44546 44942 44548 44994
rect 44492 44940 44548 44942
rect 41580 43484 41636 43540
rect 41692 43596 41748 43652
rect 41356 42812 41412 42868
rect 40236 42588 40292 42644
rect 40460 42588 40516 42644
rect 36988 42364 37044 42420
rect 37772 41916 37828 41972
rect 39900 41858 39956 41860
rect 39900 41806 39902 41858
rect 39902 41806 39954 41858
rect 39954 41806 39956 41858
rect 39900 41804 39956 41806
rect 44044 42866 44100 42868
rect 44044 42814 44046 42866
rect 44046 42814 44098 42866
rect 44098 42814 44100 42866
rect 44044 42812 44100 42814
rect 41916 42642 41972 42644
rect 41916 42590 41918 42642
rect 41918 42590 41970 42642
rect 41970 42590 41972 42642
rect 41916 42588 41972 42590
rect 44828 52834 44884 52836
rect 44828 52782 44830 52834
rect 44830 52782 44882 52834
rect 44882 52782 44884 52834
rect 44828 52780 44884 52782
rect 45388 48860 45444 48916
rect 54460 56252 54516 56308
rect 56028 56306 56084 56308
rect 56028 56254 56030 56306
rect 56030 56254 56082 56306
rect 56082 56254 56084 56306
rect 56028 56252 56084 56254
rect 52332 55356 52388 55412
rect 53676 55410 53732 55412
rect 53676 55358 53678 55410
rect 53678 55358 53730 55410
rect 53730 55358 53732 55410
rect 53676 55356 53732 55358
rect 50556 54906 50612 54908
rect 50556 54854 50558 54906
rect 50558 54854 50610 54906
rect 50610 54854 50612 54906
rect 50556 54852 50612 54854
rect 50660 54906 50716 54908
rect 50660 54854 50662 54906
rect 50662 54854 50714 54906
rect 50714 54854 50716 54906
rect 50660 54852 50716 54854
rect 50764 54906 50820 54908
rect 50764 54854 50766 54906
rect 50766 54854 50818 54906
rect 50818 54854 50820 54906
rect 50764 54852 50820 54854
rect 47740 47516 47796 47572
rect 50556 53338 50612 53340
rect 50556 53286 50558 53338
rect 50558 53286 50610 53338
rect 50610 53286 50612 53338
rect 50556 53284 50612 53286
rect 50660 53338 50716 53340
rect 50660 53286 50662 53338
rect 50662 53286 50714 53338
rect 50714 53286 50716 53338
rect 50660 53284 50716 53286
rect 50764 53338 50820 53340
rect 50764 53286 50766 53338
rect 50766 53286 50818 53338
rect 50818 53286 50820 53338
rect 50764 53284 50820 53286
rect 50556 51770 50612 51772
rect 50556 51718 50558 51770
rect 50558 51718 50610 51770
rect 50610 51718 50612 51770
rect 50556 51716 50612 51718
rect 50660 51770 50716 51772
rect 50660 51718 50662 51770
rect 50662 51718 50714 51770
rect 50714 51718 50716 51770
rect 50660 51716 50716 51718
rect 50764 51770 50820 51772
rect 50764 51718 50766 51770
rect 50766 51718 50818 51770
rect 50818 51718 50820 51770
rect 50764 51716 50820 51718
rect 50556 50202 50612 50204
rect 50556 50150 50558 50202
rect 50558 50150 50610 50202
rect 50610 50150 50612 50202
rect 50556 50148 50612 50150
rect 50660 50202 50716 50204
rect 50660 50150 50662 50202
rect 50662 50150 50714 50202
rect 50714 50150 50716 50202
rect 50660 50148 50716 50150
rect 50764 50202 50820 50204
rect 50764 50150 50766 50202
rect 50766 50150 50818 50202
rect 50818 50150 50820 50202
rect 50764 50148 50820 50150
rect 50556 48634 50612 48636
rect 50556 48582 50558 48634
rect 50558 48582 50610 48634
rect 50610 48582 50612 48634
rect 50556 48580 50612 48582
rect 50660 48634 50716 48636
rect 50660 48582 50662 48634
rect 50662 48582 50714 48634
rect 50714 48582 50716 48634
rect 50660 48580 50716 48582
rect 50764 48634 50820 48636
rect 50764 48582 50766 48634
rect 50766 48582 50818 48634
rect 50818 48582 50820 48634
rect 50764 48580 50820 48582
rect 50556 47066 50612 47068
rect 50556 47014 50558 47066
rect 50558 47014 50610 47066
rect 50610 47014 50612 47066
rect 50556 47012 50612 47014
rect 50660 47066 50716 47068
rect 50660 47014 50662 47066
rect 50662 47014 50714 47066
rect 50714 47014 50716 47066
rect 50660 47012 50716 47014
rect 50764 47066 50820 47068
rect 50764 47014 50766 47066
rect 50766 47014 50818 47066
rect 50818 47014 50820 47066
rect 50764 47012 50820 47014
rect 50316 45948 50372 46004
rect 50556 45498 50612 45500
rect 50556 45446 50558 45498
rect 50558 45446 50610 45498
rect 50610 45446 50612 45498
rect 50556 45444 50612 45446
rect 50660 45498 50716 45500
rect 50660 45446 50662 45498
rect 50662 45446 50714 45498
rect 50714 45446 50716 45498
rect 50660 45444 50716 45446
rect 50764 45498 50820 45500
rect 50764 45446 50766 45498
rect 50766 45446 50818 45498
rect 50818 45446 50820 45498
rect 50764 45444 50820 45446
rect 50556 43930 50612 43932
rect 50556 43878 50558 43930
rect 50558 43878 50610 43930
rect 50610 43878 50612 43930
rect 50556 43876 50612 43878
rect 50660 43930 50716 43932
rect 50660 43878 50662 43930
rect 50662 43878 50714 43930
rect 50714 43878 50716 43930
rect 50660 43876 50716 43878
rect 50764 43930 50820 43932
rect 50764 43878 50766 43930
rect 50766 43878 50818 43930
rect 50818 43878 50820 43930
rect 50764 43876 50820 43878
rect 44604 42364 44660 42420
rect 50556 42362 50612 42364
rect 50556 42310 50558 42362
rect 50558 42310 50610 42362
rect 50610 42310 50612 42362
rect 50556 42308 50612 42310
rect 50660 42362 50716 42364
rect 50660 42310 50662 42362
rect 50662 42310 50714 42362
rect 50714 42310 50716 42362
rect 50660 42308 50716 42310
rect 50764 42362 50820 42364
rect 50764 42310 50766 42362
rect 50766 42310 50818 42362
rect 50818 42310 50820 42362
rect 50764 42308 50820 42310
rect 40460 41804 40516 41860
rect 40908 41132 40964 41188
rect 54572 53788 54628 53844
rect 55356 44380 55412 44436
rect 52108 40908 52164 40964
rect 50556 40794 50612 40796
rect 50556 40742 50558 40794
rect 50558 40742 50610 40794
rect 50610 40742 50612 40794
rect 50556 40740 50612 40742
rect 50660 40794 50716 40796
rect 50660 40742 50662 40794
rect 50662 40742 50714 40794
rect 50714 40742 50716 40794
rect 50660 40740 50716 40742
rect 50764 40794 50820 40796
rect 50764 40742 50766 40794
rect 50766 40742 50818 40794
rect 50818 40742 50820 40794
rect 50764 40740 50820 40742
rect 36428 37996 36484 38052
rect 35644 37212 35700 37268
rect 38220 38946 38276 38948
rect 38220 38894 38222 38946
rect 38222 38894 38274 38946
rect 38274 38894 38276 38946
rect 38220 38892 38276 38894
rect 36988 38668 37044 38724
rect 37436 38668 37492 38724
rect 37212 38220 37268 38276
rect 37772 38274 37828 38276
rect 37772 38222 37774 38274
rect 37774 38222 37826 38274
rect 37826 38222 37828 38274
rect 37772 38220 37828 38222
rect 50556 39226 50612 39228
rect 50556 39174 50558 39226
rect 50558 39174 50610 39226
rect 50610 39174 50612 39226
rect 50556 39172 50612 39174
rect 50660 39226 50716 39228
rect 50660 39174 50662 39226
rect 50662 39174 50714 39226
rect 50714 39174 50716 39226
rect 50660 39172 50716 39174
rect 50764 39226 50820 39228
rect 50764 39174 50766 39226
rect 50766 39174 50818 39226
rect 50818 39174 50820 39226
rect 50764 39172 50820 39174
rect 39340 38220 39396 38276
rect 37996 37154 38052 37156
rect 37996 37102 37998 37154
rect 37998 37102 38050 37154
rect 38050 37102 38052 37154
rect 37996 37100 38052 37102
rect 38444 38050 38500 38052
rect 38444 37998 38446 38050
rect 38446 37998 38498 38050
rect 38498 37998 38500 38050
rect 38444 37996 38500 37998
rect 38108 37324 38164 37380
rect 35532 35868 35588 35924
rect 35644 35756 35700 35812
rect 34748 35420 34804 35476
rect 34972 35698 35028 35700
rect 34972 35646 34974 35698
rect 34974 35646 35026 35698
rect 35026 35646 35028 35698
rect 34972 35644 35028 35646
rect 34524 32620 34580 32676
rect 34748 32844 34804 32900
rect 34748 32508 34804 32564
rect 34412 31052 34468 31108
rect 35196 35306 35252 35308
rect 35196 35254 35198 35306
rect 35198 35254 35250 35306
rect 35250 35254 35252 35306
rect 35196 35252 35252 35254
rect 35300 35306 35356 35308
rect 35300 35254 35302 35306
rect 35302 35254 35354 35306
rect 35354 35254 35356 35306
rect 35300 35252 35356 35254
rect 35404 35306 35460 35308
rect 35404 35254 35406 35306
rect 35406 35254 35458 35306
rect 35458 35254 35460 35306
rect 35404 35252 35460 35254
rect 36428 35868 36484 35924
rect 36204 35644 36260 35700
rect 37100 35698 37156 35700
rect 37100 35646 37102 35698
rect 37102 35646 37154 35698
rect 37154 35646 37156 35698
rect 37100 35644 37156 35646
rect 35532 35084 35588 35140
rect 35308 34690 35364 34692
rect 35308 34638 35310 34690
rect 35310 34638 35362 34690
rect 35362 34638 35364 34690
rect 35308 34636 35364 34638
rect 36316 35420 36372 35476
rect 36316 34802 36372 34804
rect 36316 34750 36318 34802
rect 36318 34750 36370 34802
rect 36370 34750 36372 34802
rect 36316 34748 36372 34750
rect 36428 35308 36484 35364
rect 36876 34860 36932 34916
rect 35420 34076 35476 34132
rect 36092 34130 36148 34132
rect 36092 34078 36094 34130
rect 36094 34078 36146 34130
rect 36146 34078 36148 34130
rect 36092 34076 36148 34078
rect 35196 33738 35252 33740
rect 35196 33686 35198 33738
rect 35198 33686 35250 33738
rect 35250 33686 35252 33738
rect 35196 33684 35252 33686
rect 35300 33738 35356 33740
rect 35300 33686 35302 33738
rect 35302 33686 35354 33738
rect 35354 33686 35356 33738
rect 35300 33684 35356 33686
rect 35404 33738 35460 33740
rect 35404 33686 35406 33738
rect 35406 33686 35458 33738
rect 35458 33686 35460 33738
rect 35404 33684 35460 33686
rect 36092 33628 36148 33684
rect 34972 32844 35028 32900
rect 36428 34130 36484 34132
rect 36428 34078 36430 34130
rect 36430 34078 36482 34130
rect 36482 34078 36484 34130
rect 36428 34076 36484 34078
rect 35196 32562 35252 32564
rect 35196 32510 35198 32562
rect 35198 32510 35250 32562
rect 35250 32510 35252 32562
rect 35196 32508 35252 32510
rect 35644 33180 35700 33236
rect 36428 32844 36484 32900
rect 35196 32170 35252 32172
rect 35196 32118 35198 32170
rect 35198 32118 35250 32170
rect 35250 32118 35252 32170
rect 35196 32116 35252 32118
rect 35300 32170 35356 32172
rect 35300 32118 35302 32170
rect 35302 32118 35354 32170
rect 35354 32118 35356 32170
rect 35300 32116 35356 32118
rect 35404 32170 35460 32172
rect 35404 32118 35406 32170
rect 35406 32118 35458 32170
rect 35458 32118 35460 32170
rect 35404 32116 35460 32118
rect 35196 31666 35252 31668
rect 35196 31614 35198 31666
rect 35198 31614 35250 31666
rect 35250 31614 35252 31666
rect 35196 31612 35252 31614
rect 35644 31612 35700 31668
rect 35756 31106 35812 31108
rect 35756 31054 35758 31106
rect 35758 31054 35810 31106
rect 35810 31054 35812 31106
rect 35756 31052 35812 31054
rect 35980 30940 36036 30996
rect 35196 30602 35252 30604
rect 35196 30550 35198 30602
rect 35198 30550 35250 30602
rect 35250 30550 35252 30602
rect 35196 30548 35252 30550
rect 35300 30602 35356 30604
rect 35300 30550 35302 30602
rect 35302 30550 35354 30602
rect 35354 30550 35356 30602
rect 35300 30548 35356 30550
rect 35404 30602 35460 30604
rect 35404 30550 35406 30602
rect 35406 30550 35458 30602
rect 35458 30550 35460 30602
rect 35404 30548 35460 30550
rect 34972 30210 35028 30212
rect 34972 30158 34974 30210
rect 34974 30158 35026 30210
rect 35026 30158 35028 30210
rect 34972 30156 35028 30158
rect 35644 30210 35700 30212
rect 35644 30158 35646 30210
rect 35646 30158 35698 30210
rect 35698 30158 35700 30210
rect 35644 30156 35700 30158
rect 35196 29034 35252 29036
rect 35196 28982 35198 29034
rect 35198 28982 35250 29034
rect 35250 28982 35252 29034
rect 35196 28980 35252 28982
rect 35300 29034 35356 29036
rect 35300 28982 35302 29034
rect 35302 28982 35354 29034
rect 35354 28982 35356 29034
rect 35300 28980 35356 28982
rect 35404 29034 35460 29036
rect 35404 28982 35406 29034
rect 35406 28982 35458 29034
rect 35458 28982 35460 29034
rect 35404 28980 35460 28982
rect 37100 34802 37156 34804
rect 37100 34750 37102 34802
rect 37102 34750 37154 34802
rect 37154 34750 37156 34802
rect 37100 34748 37156 34750
rect 37212 34690 37268 34692
rect 37212 34638 37214 34690
rect 37214 34638 37266 34690
rect 37266 34638 37268 34690
rect 37212 34636 37268 34638
rect 37996 36482 38052 36484
rect 37996 36430 37998 36482
rect 37998 36430 38050 36482
rect 38050 36430 38052 36482
rect 37996 36428 38052 36430
rect 38668 37100 38724 37156
rect 38444 35980 38500 36036
rect 37436 35810 37492 35812
rect 37436 35758 37438 35810
rect 37438 35758 37490 35810
rect 37490 35758 37492 35810
rect 37436 35756 37492 35758
rect 37660 34748 37716 34804
rect 37324 33628 37380 33684
rect 37100 33346 37156 33348
rect 37100 33294 37102 33346
rect 37102 33294 37154 33346
rect 37154 33294 37156 33346
rect 37100 33292 37156 33294
rect 37212 33122 37268 33124
rect 37212 33070 37214 33122
rect 37214 33070 37266 33122
rect 37266 33070 37268 33122
rect 37212 33068 37268 33070
rect 37660 32732 37716 32788
rect 37324 32674 37380 32676
rect 37324 32622 37326 32674
rect 37326 32622 37378 32674
rect 37378 32622 37380 32674
rect 37324 32620 37380 32622
rect 36876 30994 36932 30996
rect 36876 30942 36878 30994
rect 36878 30942 36930 30994
rect 36930 30942 36932 30994
rect 36876 30940 36932 30942
rect 35980 30098 36036 30100
rect 35980 30046 35982 30098
rect 35982 30046 36034 30098
rect 36034 30046 36036 30098
rect 35980 30044 36036 30046
rect 35756 28028 35812 28084
rect 35196 27466 35252 27468
rect 35196 27414 35198 27466
rect 35198 27414 35250 27466
rect 35250 27414 35252 27466
rect 35196 27412 35252 27414
rect 35300 27466 35356 27468
rect 35300 27414 35302 27466
rect 35302 27414 35354 27466
rect 35354 27414 35356 27466
rect 35300 27412 35356 27414
rect 35404 27466 35460 27468
rect 35404 27414 35406 27466
rect 35406 27414 35458 27466
rect 35458 27414 35460 27466
rect 35404 27412 35460 27414
rect 28252 26572 28308 26628
rect 29260 25282 29316 25284
rect 29260 25230 29262 25282
rect 29262 25230 29314 25282
rect 29314 25230 29316 25282
rect 29260 25228 29316 25230
rect 35196 25898 35252 25900
rect 35196 25846 35198 25898
rect 35198 25846 35250 25898
rect 35250 25846 35252 25898
rect 35196 25844 35252 25846
rect 35300 25898 35356 25900
rect 35300 25846 35302 25898
rect 35302 25846 35354 25898
rect 35354 25846 35356 25898
rect 35300 25844 35356 25846
rect 35404 25898 35460 25900
rect 35404 25846 35406 25898
rect 35406 25846 35458 25898
rect 35458 25846 35460 25898
rect 35404 25844 35460 25846
rect 33628 25564 33684 25620
rect 37436 31612 37492 31668
rect 37212 31554 37268 31556
rect 37212 31502 37214 31554
rect 37214 31502 37266 31554
rect 37266 31502 37268 31554
rect 37212 31500 37268 31502
rect 36988 30156 37044 30212
rect 37212 30210 37268 30212
rect 37212 30158 37214 30210
rect 37214 30158 37266 30210
rect 37266 30158 37268 30210
rect 37212 30156 37268 30158
rect 36540 30098 36596 30100
rect 36540 30046 36542 30098
rect 36542 30046 36594 30098
rect 36594 30046 36596 30098
rect 36540 30044 36596 30046
rect 39004 36204 39060 36260
rect 39004 35644 39060 35700
rect 38668 35084 38724 35140
rect 38556 34914 38612 34916
rect 38556 34862 38558 34914
rect 38558 34862 38610 34914
rect 38610 34862 38612 34914
rect 38556 34860 38612 34862
rect 39228 35868 39284 35924
rect 39116 35308 39172 35364
rect 38220 33628 38276 33684
rect 38892 33628 38948 33684
rect 39340 35084 39396 35140
rect 39900 38220 39956 38276
rect 50556 37658 50612 37660
rect 50556 37606 50558 37658
rect 50558 37606 50610 37658
rect 50610 37606 50612 37658
rect 50556 37604 50612 37606
rect 50660 37658 50716 37660
rect 50660 37606 50662 37658
rect 50662 37606 50714 37658
rect 50714 37606 50716 37658
rect 50660 37604 50716 37606
rect 50764 37658 50820 37660
rect 50764 37606 50766 37658
rect 50766 37606 50818 37658
rect 50818 37606 50820 37658
rect 50764 37604 50820 37606
rect 39564 37378 39620 37380
rect 39564 37326 39566 37378
rect 39566 37326 39618 37378
rect 39618 37326 39620 37378
rect 39564 37324 39620 37326
rect 40124 36258 40180 36260
rect 40124 36206 40126 36258
rect 40126 36206 40178 36258
rect 40178 36206 40180 36258
rect 40124 36204 40180 36206
rect 40348 35980 40404 36036
rect 40908 35980 40964 36036
rect 39676 35532 39732 35588
rect 39564 34076 39620 34132
rect 40124 34076 40180 34132
rect 39452 33292 39508 33348
rect 39676 33516 39732 33572
rect 38668 33068 38724 33124
rect 39116 32844 39172 32900
rect 38108 30156 38164 30212
rect 40908 33292 40964 33348
rect 50556 36090 50612 36092
rect 50556 36038 50558 36090
rect 50558 36038 50610 36090
rect 50610 36038 50612 36090
rect 50556 36036 50612 36038
rect 50660 36090 50716 36092
rect 50660 36038 50662 36090
rect 50662 36038 50714 36090
rect 50714 36038 50716 36090
rect 50660 36036 50716 36038
rect 50764 36090 50820 36092
rect 50764 36038 50766 36090
rect 50766 36038 50818 36090
rect 50818 36038 50820 36090
rect 50764 36036 50820 36038
rect 41356 35586 41412 35588
rect 41356 35534 41358 35586
rect 41358 35534 41410 35586
rect 41410 35534 41412 35586
rect 41356 35532 41412 35534
rect 41468 34748 41524 34804
rect 50556 34522 50612 34524
rect 50556 34470 50558 34522
rect 50558 34470 50610 34522
rect 50610 34470 50612 34522
rect 50556 34468 50612 34470
rect 50660 34522 50716 34524
rect 50660 34470 50662 34522
rect 50662 34470 50714 34522
rect 50714 34470 50716 34522
rect 50660 34468 50716 34470
rect 50764 34522 50820 34524
rect 50764 34470 50766 34522
rect 50766 34470 50818 34522
rect 50818 34470 50820 34522
rect 50764 34468 50820 34470
rect 50556 32954 50612 32956
rect 50556 32902 50558 32954
rect 50558 32902 50610 32954
rect 50610 32902 50612 32954
rect 50556 32900 50612 32902
rect 50660 32954 50716 32956
rect 50660 32902 50662 32954
rect 50662 32902 50714 32954
rect 50714 32902 50716 32954
rect 50660 32900 50716 32902
rect 50764 32954 50820 32956
rect 50764 32902 50766 32954
rect 50766 32902 50818 32954
rect 50818 32902 50820 32954
rect 50764 32900 50820 32902
rect 50556 31386 50612 31388
rect 50556 31334 50558 31386
rect 50558 31334 50610 31386
rect 50610 31334 50612 31386
rect 50556 31332 50612 31334
rect 50660 31386 50716 31388
rect 50660 31334 50662 31386
rect 50662 31334 50714 31386
rect 50714 31334 50716 31386
rect 50660 31332 50716 31334
rect 50764 31386 50820 31388
rect 50764 31334 50766 31386
rect 50766 31334 50818 31386
rect 50818 31334 50820 31386
rect 50764 31332 50820 31334
rect 39452 31052 39508 31108
rect 50556 29818 50612 29820
rect 50556 29766 50558 29818
rect 50558 29766 50610 29818
rect 50610 29766 50612 29818
rect 50556 29764 50612 29766
rect 50660 29818 50716 29820
rect 50660 29766 50662 29818
rect 50662 29766 50714 29818
rect 50714 29766 50716 29818
rect 50660 29764 50716 29766
rect 50764 29818 50820 29820
rect 50764 29766 50766 29818
rect 50766 29766 50818 29818
rect 50818 29766 50820 29818
rect 50764 29764 50820 29766
rect 50556 28250 50612 28252
rect 50556 28198 50558 28250
rect 50558 28198 50610 28250
rect 50610 28198 50612 28250
rect 50556 28196 50612 28198
rect 50660 28250 50716 28252
rect 50660 28198 50662 28250
rect 50662 28198 50714 28250
rect 50714 28198 50716 28250
rect 50660 28196 50716 28198
rect 50764 28250 50820 28252
rect 50764 28198 50766 28250
rect 50766 28198 50818 28250
rect 50818 28198 50820 28250
rect 50764 28196 50820 28198
rect 50556 26682 50612 26684
rect 50556 26630 50558 26682
rect 50558 26630 50610 26682
rect 50610 26630 50612 26682
rect 50556 26628 50612 26630
rect 50660 26682 50716 26684
rect 50660 26630 50662 26682
rect 50662 26630 50714 26682
rect 50714 26630 50716 26682
rect 50660 26628 50716 26630
rect 50764 26682 50820 26684
rect 50764 26630 50766 26682
rect 50766 26630 50818 26682
rect 50818 26630 50820 26682
rect 50764 26628 50820 26630
rect 36428 25228 36484 25284
rect 50556 25114 50612 25116
rect 50556 25062 50558 25114
rect 50558 25062 50610 25114
rect 50610 25062 50612 25114
rect 50556 25060 50612 25062
rect 50660 25114 50716 25116
rect 50660 25062 50662 25114
rect 50662 25062 50714 25114
rect 50714 25062 50716 25114
rect 50660 25060 50716 25062
rect 50764 25114 50820 25116
rect 50764 25062 50766 25114
rect 50766 25062 50818 25114
rect 50818 25062 50820 25114
rect 50764 25060 50820 25062
rect 32060 24892 32116 24948
rect 30492 24780 30548 24836
rect 35196 24330 35252 24332
rect 35196 24278 35198 24330
rect 35198 24278 35250 24330
rect 35250 24278 35252 24330
rect 35196 24276 35252 24278
rect 35300 24330 35356 24332
rect 35300 24278 35302 24330
rect 35302 24278 35354 24330
rect 35354 24278 35356 24330
rect 35300 24276 35356 24278
rect 35404 24330 35460 24332
rect 35404 24278 35406 24330
rect 35406 24278 35458 24330
rect 35458 24278 35460 24330
rect 35404 24276 35460 24278
rect 50556 23546 50612 23548
rect 50556 23494 50558 23546
rect 50558 23494 50610 23546
rect 50610 23494 50612 23546
rect 50556 23492 50612 23494
rect 50660 23546 50716 23548
rect 50660 23494 50662 23546
rect 50662 23494 50714 23546
rect 50714 23494 50716 23546
rect 50660 23492 50716 23494
rect 50764 23546 50820 23548
rect 50764 23494 50766 23546
rect 50766 23494 50818 23546
rect 50818 23494 50820 23546
rect 50764 23492 50820 23494
rect 27916 22876 27972 22932
rect 27804 22652 27860 22708
rect 35196 22762 35252 22764
rect 35196 22710 35198 22762
rect 35198 22710 35250 22762
rect 35250 22710 35252 22762
rect 35196 22708 35252 22710
rect 35300 22762 35356 22764
rect 35300 22710 35302 22762
rect 35302 22710 35354 22762
rect 35354 22710 35356 22762
rect 35300 22708 35356 22710
rect 35404 22762 35460 22764
rect 35404 22710 35406 22762
rect 35406 22710 35458 22762
rect 35458 22710 35460 22762
rect 35404 22708 35460 22710
rect 19836 21978 19892 21980
rect 19836 21926 19838 21978
rect 19838 21926 19890 21978
rect 19890 21926 19892 21978
rect 19836 21924 19892 21926
rect 19940 21978 19996 21980
rect 19940 21926 19942 21978
rect 19942 21926 19994 21978
rect 19994 21926 19996 21978
rect 19940 21924 19996 21926
rect 20044 21978 20100 21980
rect 20044 21926 20046 21978
rect 20046 21926 20098 21978
rect 20098 21926 20100 21978
rect 20044 21924 20100 21926
rect 50556 21978 50612 21980
rect 50556 21926 50558 21978
rect 50558 21926 50610 21978
rect 50610 21926 50612 21978
rect 50556 21924 50612 21926
rect 50660 21978 50716 21980
rect 50660 21926 50662 21978
rect 50662 21926 50714 21978
rect 50714 21926 50716 21978
rect 50660 21924 50716 21926
rect 50764 21978 50820 21980
rect 50764 21926 50766 21978
rect 50766 21926 50818 21978
rect 50818 21926 50820 21978
rect 50764 21924 50820 21926
rect 12684 21644 12740 21700
rect 35196 21194 35252 21196
rect 35196 21142 35198 21194
rect 35198 21142 35250 21194
rect 35250 21142 35252 21194
rect 35196 21140 35252 21142
rect 35300 21194 35356 21196
rect 35300 21142 35302 21194
rect 35302 21142 35354 21194
rect 35354 21142 35356 21194
rect 35300 21140 35356 21142
rect 35404 21194 35460 21196
rect 35404 21142 35406 21194
rect 35406 21142 35458 21194
rect 35458 21142 35460 21194
rect 35404 21140 35460 21142
rect 19836 20410 19892 20412
rect 19836 20358 19838 20410
rect 19838 20358 19890 20410
rect 19890 20358 19892 20410
rect 19836 20356 19892 20358
rect 19940 20410 19996 20412
rect 19940 20358 19942 20410
rect 19942 20358 19994 20410
rect 19994 20358 19996 20410
rect 19940 20356 19996 20358
rect 20044 20410 20100 20412
rect 20044 20358 20046 20410
rect 20046 20358 20098 20410
rect 20098 20358 20100 20410
rect 20044 20356 20100 20358
rect 50556 20410 50612 20412
rect 50556 20358 50558 20410
rect 50558 20358 50610 20410
rect 50610 20358 50612 20410
rect 50556 20356 50612 20358
rect 50660 20410 50716 20412
rect 50660 20358 50662 20410
rect 50662 20358 50714 20410
rect 50714 20358 50716 20410
rect 50660 20356 50716 20358
rect 50764 20410 50820 20412
rect 50764 20358 50766 20410
rect 50766 20358 50818 20410
rect 50818 20358 50820 20410
rect 50764 20356 50820 20358
rect 6524 9996 6580 10052
rect 2492 9212 2548 9268
rect 4476 8650 4532 8652
rect 4476 8598 4478 8650
rect 4478 8598 4530 8650
rect 4530 8598 4532 8650
rect 4476 8596 4532 8598
rect 4580 8650 4636 8652
rect 4580 8598 4582 8650
rect 4582 8598 4634 8650
rect 4634 8598 4636 8650
rect 4580 8596 4636 8598
rect 4684 8650 4740 8652
rect 4684 8598 4686 8650
rect 4686 8598 4738 8650
rect 4738 8598 4740 8650
rect 4684 8596 4740 8598
rect 2492 8034 2548 8036
rect 2492 7982 2494 8034
rect 2494 7982 2546 8034
rect 2546 7982 2548 8034
rect 2492 7980 2548 7982
rect 4476 7082 4532 7084
rect 4476 7030 4478 7082
rect 4478 7030 4530 7082
rect 4530 7030 4532 7082
rect 4476 7028 4532 7030
rect 4580 7082 4636 7084
rect 4580 7030 4582 7082
rect 4582 7030 4634 7082
rect 4634 7030 4636 7082
rect 4580 7028 4636 7030
rect 4684 7082 4740 7084
rect 4684 7030 4686 7082
rect 4686 7030 4738 7082
rect 4738 7030 4740 7082
rect 4684 7028 4740 7030
rect 4476 5514 4532 5516
rect 4476 5462 4478 5514
rect 4478 5462 4530 5514
rect 4530 5462 4532 5514
rect 4476 5460 4532 5462
rect 4580 5514 4636 5516
rect 4580 5462 4582 5514
rect 4582 5462 4634 5514
rect 4634 5462 4636 5514
rect 4580 5460 4636 5462
rect 4684 5514 4740 5516
rect 4684 5462 4686 5514
rect 4686 5462 4738 5514
rect 4738 5462 4740 5514
rect 4684 5460 4740 5462
rect 35196 19626 35252 19628
rect 35196 19574 35198 19626
rect 35198 19574 35250 19626
rect 35250 19574 35252 19626
rect 35196 19572 35252 19574
rect 35300 19626 35356 19628
rect 35300 19574 35302 19626
rect 35302 19574 35354 19626
rect 35354 19574 35356 19626
rect 35300 19572 35356 19574
rect 35404 19626 35460 19628
rect 35404 19574 35406 19626
rect 35406 19574 35458 19626
rect 35458 19574 35460 19626
rect 35404 19572 35460 19574
rect 19836 18842 19892 18844
rect 19836 18790 19838 18842
rect 19838 18790 19890 18842
rect 19890 18790 19892 18842
rect 19836 18788 19892 18790
rect 19940 18842 19996 18844
rect 19940 18790 19942 18842
rect 19942 18790 19994 18842
rect 19994 18790 19996 18842
rect 19940 18788 19996 18790
rect 20044 18842 20100 18844
rect 20044 18790 20046 18842
rect 20046 18790 20098 18842
rect 20098 18790 20100 18842
rect 20044 18788 20100 18790
rect 50556 18842 50612 18844
rect 50556 18790 50558 18842
rect 50558 18790 50610 18842
rect 50610 18790 50612 18842
rect 50556 18788 50612 18790
rect 50660 18842 50716 18844
rect 50660 18790 50662 18842
rect 50662 18790 50714 18842
rect 50714 18790 50716 18842
rect 50660 18788 50716 18790
rect 50764 18842 50820 18844
rect 50764 18790 50766 18842
rect 50766 18790 50818 18842
rect 50818 18790 50820 18842
rect 50764 18788 50820 18790
rect 35196 18058 35252 18060
rect 35196 18006 35198 18058
rect 35198 18006 35250 18058
rect 35250 18006 35252 18058
rect 35196 18004 35252 18006
rect 35300 18058 35356 18060
rect 35300 18006 35302 18058
rect 35302 18006 35354 18058
rect 35354 18006 35356 18058
rect 35300 18004 35356 18006
rect 35404 18058 35460 18060
rect 35404 18006 35406 18058
rect 35406 18006 35458 18058
rect 35458 18006 35460 18058
rect 35404 18004 35460 18006
rect 19836 17274 19892 17276
rect 19836 17222 19838 17274
rect 19838 17222 19890 17274
rect 19890 17222 19892 17274
rect 19836 17220 19892 17222
rect 19940 17274 19996 17276
rect 19940 17222 19942 17274
rect 19942 17222 19994 17274
rect 19994 17222 19996 17274
rect 19940 17220 19996 17222
rect 20044 17274 20100 17276
rect 20044 17222 20046 17274
rect 20046 17222 20098 17274
rect 20098 17222 20100 17274
rect 20044 17220 20100 17222
rect 50556 17274 50612 17276
rect 50556 17222 50558 17274
rect 50558 17222 50610 17274
rect 50610 17222 50612 17274
rect 50556 17220 50612 17222
rect 50660 17274 50716 17276
rect 50660 17222 50662 17274
rect 50662 17222 50714 17274
rect 50714 17222 50716 17274
rect 50660 17220 50716 17222
rect 50764 17274 50820 17276
rect 50764 17222 50766 17274
rect 50766 17222 50818 17274
rect 50818 17222 50820 17274
rect 50764 17220 50820 17222
rect 35196 16490 35252 16492
rect 35196 16438 35198 16490
rect 35198 16438 35250 16490
rect 35250 16438 35252 16490
rect 35196 16436 35252 16438
rect 35300 16490 35356 16492
rect 35300 16438 35302 16490
rect 35302 16438 35354 16490
rect 35354 16438 35356 16490
rect 35300 16436 35356 16438
rect 35404 16490 35460 16492
rect 35404 16438 35406 16490
rect 35406 16438 35458 16490
rect 35458 16438 35460 16490
rect 35404 16436 35460 16438
rect 19836 15706 19892 15708
rect 19836 15654 19838 15706
rect 19838 15654 19890 15706
rect 19890 15654 19892 15706
rect 19836 15652 19892 15654
rect 19940 15706 19996 15708
rect 19940 15654 19942 15706
rect 19942 15654 19994 15706
rect 19994 15654 19996 15706
rect 19940 15652 19996 15654
rect 20044 15706 20100 15708
rect 20044 15654 20046 15706
rect 20046 15654 20098 15706
rect 20098 15654 20100 15706
rect 20044 15652 20100 15654
rect 50556 15706 50612 15708
rect 50556 15654 50558 15706
rect 50558 15654 50610 15706
rect 50610 15654 50612 15706
rect 50556 15652 50612 15654
rect 50660 15706 50716 15708
rect 50660 15654 50662 15706
rect 50662 15654 50714 15706
rect 50714 15654 50716 15706
rect 50660 15652 50716 15654
rect 50764 15706 50820 15708
rect 50764 15654 50766 15706
rect 50766 15654 50818 15706
rect 50818 15654 50820 15706
rect 50764 15652 50820 15654
rect 35196 14922 35252 14924
rect 35196 14870 35198 14922
rect 35198 14870 35250 14922
rect 35250 14870 35252 14922
rect 35196 14868 35252 14870
rect 35300 14922 35356 14924
rect 35300 14870 35302 14922
rect 35302 14870 35354 14922
rect 35354 14870 35356 14922
rect 35300 14868 35356 14870
rect 35404 14922 35460 14924
rect 35404 14870 35406 14922
rect 35406 14870 35458 14922
rect 35458 14870 35460 14922
rect 35404 14868 35460 14870
rect 19836 14138 19892 14140
rect 19836 14086 19838 14138
rect 19838 14086 19890 14138
rect 19890 14086 19892 14138
rect 19836 14084 19892 14086
rect 19940 14138 19996 14140
rect 19940 14086 19942 14138
rect 19942 14086 19994 14138
rect 19994 14086 19996 14138
rect 19940 14084 19996 14086
rect 20044 14138 20100 14140
rect 20044 14086 20046 14138
rect 20046 14086 20098 14138
rect 20098 14086 20100 14138
rect 20044 14084 20100 14086
rect 50556 14138 50612 14140
rect 50556 14086 50558 14138
rect 50558 14086 50610 14138
rect 50610 14086 50612 14138
rect 50556 14084 50612 14086
rect 50660 14138 50716 14140
rect 50660 14086 50662 14138
rect 50662 14086 50714 14138
rect 50714 14086 50716 14138
rect 50660 14084 50716 14086
rect 50764 14138 50820 14140
rect 50764 14086 50766 14138
rect 50766 14086 50818 14138
rect 50818 14086 50820 14138
rect 50764 14084 50820 14086
rect 35196 13354 35252 13356
rect 35196 13302 35198 13354
rect 35198 13302 35250 13354
rect 35250 13302 35252 13354
rect 35196 13300 35252 13302
rect 35300 13354 35356 13356
rect 35300 13302 35302 13354
rect 35302 13302 35354 13354
rect 35354 13302 35356 13354
rect 35300 13300 35356 13302
rect 35404 13354 35460 13356
rect 35404 13302 35406 13354
rect 35406 13302 35458 13354
rect 35458 13302 35460 13354
rect 35404 13300 35460 13302
rect 19836 12570 19892 12572
rect 19836 12518 19838 12570
rect 19838 12518 19890 12570
rect 19890 12518 19892 12570
rect 19836 12516 19892 12518
rect 19940 12570 19996 12572
rect 19940 12518 19942 12570
rect 19942 12518 19994 12570
rect 19994 12518 19996 12570
rect 19940 12516 19996 12518
rect 20044 12570 20100 12572
rect 20044 12518 20046 12570
rect 20046 12518 20098 12570
rect 20098 12518 20100 12570
rect 20044 12516 20100 12518
rect 50556 12570 50612 12572
rect 50556 12518 50558 12570
rect 50558 12518 50610 12570
rect 50610 12518 50612 12570
rect 50556 12516 50612 12518
rect 50660 12570 50716 12572
rect 50660 12518 50662 12570
rect 50662 12518 50714 12570
rect 50714 12518 50716 12570
rect 50660 12516 50716 12518
rect 50764 12570 50820 12572
rect 50764 12518 50766 12570
rect 50766 12518 50818 12570
rect 50818 12518 50820 12570
rect 50764 12516 50820 12518
rect 35196 11786 35252 11788
rect 35196 11734 35198 11786
rect 35198 11734 35250 11786
rect 35250 11734 35252 11786
rect 35196 11732 35252 11734
rect 35300 11786 35356 11788
rect 35300 11734 35302 11786
rect 35302 11734 35354 11786
rect 35354 11734 35356 11786
rect 35300 11732 35356 11734
rect 35404 11786 35460 11788
rect 35404 11734 35406 11786
rect 35406 11734 35458 11786
rect 35458 11734 35460 11786
rect 35404 11732 35460 11734
rect 19836 11002 19892 11004
rect 19836 10950 19838 11002
rect 19838 10950 19890 11002
rect 19890 10950 19892 11002
rect 19836 10948 19892 10950
rect 19940 11002 19996 11004
rect 19940 10950 19942 11002
rect 19942 10950 19994 11002
rect 19994 10950 19996 11002
rect 19940 10948 19996 10950
rect 20044 11002 20100 11004
rect 20044 10950 20046 11002
rect 20046 10950 20098 11002
rect 20098 10950 20100 11002
rect 20044 10948 20100 10950
rect 50556 11002 50612 11004
rect 50556 10950 50558 11002
rect 50558 10950 50610 11002
rect 50610 10950 50612 11002
rect 50556 10948 50612 10950
rect 50660 11002 50716 11004
rect 50660 10950 50662 11002
rect 50662 10950 50714 11002
rect 50714 10950 50716 11002
rect 50660 10948 50716 10950
rect 50764 11002 50820 11004
rect 50764 10950 50766 11002
rect 50766 10950 50818 11002
rect 50818 10950 50820 11002
rect 50764 10948 50820 10950
rect 35196 10218 35252 10220
rect 35196 10166 35198 10218
rect 35198 10166 35250 10218
rect 35250 10166 35252 10218
rect 35196 10164 35252 10166
rect 35300 10218 35356 10220
rect 35300 10166 35302 10218
rect 35302 10166 35354 10218
rect 35354 10166 35356 10218
rect 35300 10164 35356 10166
rect 35404 10218 35460 10220
rect 35404 10166 35406 10218
rect 35406 10166 35458 10218
rect 35458 10166 35460 10218
rect 35404 10164 35460 10166
rect 19836 9434 19892 9436
rect 19836 9382 19838 9434
rect 19838 9382 19890 9434
rect 19890 9382 19892 9434
rect 19836 9380 19892 9382
rect 19940 9434 19996 9436
rect 19940 9382 19942 9434
rect 19942 9382 19994 9434
rect 19994 9382 19996 9434
rect 19940 9380 19996 9382
rect 20044 9434 20100 9436
rect 20044 9382 20046 9434
rect 20046 9382 20098 9434
rect 20098 9382 20100 9434
rect 20044 9380 20100 9382
rect 50556 9434 50612 9436
rect 50556 9382 50558 9434
rect 50558 9382 50610 9434
rect 50610 9382 50612 9434
rect 50556 9380 50612 9382
rect 50660 9434 50716 9436
rect 50660 9382 50662 9434
rect 50662 9382 50714 9434
rect 50714 9382 50716 9434
rect 50660 9380 50716 9382
rect 50764 9434 50820 9436
rect 50764 9382 50766 9434
rect 50766 9382 50818 9434
rect 50818 9382 50820 9434
rect 50764 9380 50820 9382
rect 35196 8650 35252 8652
rect 35196 8598 35198 8650
rect 35198 8598 35250 8650
rect 35250 8598 35252 8650
rect 35196 8596 35252 8598
rect 35300 8650 35356 8652
rect 35300 8598 35302 8650
rect 35302 8598 35354 8650
rect 35354 8598 35356 8650
rect 35300 8596 35356 8598
rect 35404 8650 35460 8652
rect 35404 8598 35406 8650
rect 35406 8598 35458 8650
rect 35458 8598 35460 8650
rect 35404 8596 35460 8598
rect 19836 7866 19892 7868
rect 19836 7814 19838 7866
rect 19838 7814 19890 7866
rect 19890 7814 19892 7866
rect 19836 7812 19892 7814
rect 19940 7866 19996 7868
rect 19940 7814 19942 7866
rect 19942 7814 19994 7866
rect 19994 7814 19996 7866
rect 19940 7812 19996 7814
rect 20044 7866 20100 7868
rect 20044 7814 20046 7866
rect 20046 7814 20098 7866
rect 20098 7814 20100 7866
rect 20044 7812 20100 7814
rect 50556 7866 50612 7868
rect 50556 7814 50558 7866
rect 50558 7814 50610 7866
rect 50610 7814 50612 7866
rect 50556 7812 50612 7814
rect 50660 7866 50716 7868
rect 50660 7814 50662 7866
rect 50662 7814 50714 7866
rect 50714 7814 50716 7866
rect 50660 7812 50716 7814
rect 50764 7866 50820 7868
rect 50764 7814 50766 7866
rect 50766 7814 50818 7866
rect 50818 7814 50820 7866
rect 50764 7812 50820 7814
rect 35196 7082 35252 7084
rect 35196 7030 35198 7082
rect 35198 7030 35250 7082
rect 35250 7030 35252 7082
rect 35196 7028 35252 7030
rect 35300 7082 35356 7084
rect 35300 7030 35302 7082
rect 35302 7030 35354 7082
rect 35354 7030 35356 7082
rect 35300 7028 35356 7030
rect 35404 7082 35460 7084
rect 35404 7030 35406 7082
rect 35406 7030 35458 7082
rect 35458 7030 35460 7082
rect 35404 7028 35460 7030
rect 19836 6298 19892 6300
rect 19836 6246 19838 6298
rect 19838 6246 19890 6298
rect 19890 6246 19892 6298
rect 19836 6244 19892 6246
rect 19940 6298 19996 6300
rect 19940 6246 19942 6298
rect 19942 6246 19994 6298
rect 19994 6246 19996 6298
rect 19940 6244 19996 6246
rect 20044 6298 20100 6300
rect 20044 6246 20046 6298
rect 20046 6246 20098 6298
rect 20098 6246 20100 6298
rect 20044 6244 20100 6246
rect 50556 6298 50612 6300
rect 50556 6246 50558 6298
rect 50558 6246 50610 6298
rect 50610 6246 50612 6298
rect 50556 6244 50612 6246
rect 50660 6298 50716 6300
rect 50660 6246 50662 6298
rect 50662 6246 50714 6298
rect 50714 6246 50716 6298
rect 50660 6244 50716 6246
rect 50764 6298 50820 6300
rect 50764 6246 50766 6298
rect 50766 6246 50818 6298
rect 50818 6246 50820 6298
rect 50764 6244 50820 6246
rect 35196 5514 35252 5516
rect 35196 5462 35198 5514
rect 35198 5462 35250 5514
rect 35250 5462 35252 5514
rect 35196 5460 35252 5462
rect 35300 5514 35356 5516
rect 35300 5462 35302 5514
rect 35302 5462 35354 5514
rect 35354 5462 35356 5514
rect 35300 5460 35356 5462
rect 35404 5514 35460 5516
rect 35404 5462 35406 5514
rect 35406 5462 35458 5514
rect 35458 5462 35460 5514
rect 35404 5460 35460 5462
rect 19836 4730 19892 4732
rect 19836 4678 19838 4730
rect 19838 4678 19890 4730
rect 19890 4678 19892 4730
rect 19836 4676 19892 4678
rect 19940 4730 19996 4732
rect 19940 4678 19942 4730
rect 19942 4678 19994 4730
rect 19994 4678 19996 4730
rect 19940 4676 19996 4678
rect 20044 4730 20100 4732
rect 20044 4678 20046 4730
rect 20046 4678 20098 4730
rect 20098 4678 20100 4730
rect 20044 4676 20100 4678
rect 50556 4730 50612 4732
rect 50556 4678 50558 4730
rect 50558 4678 50610 4730
rect 50610 4678 50612 4730
rect 50556 4676 50612 4678
rect 50660 4730 50716 4732
rect 50660 4678 50662 4730
rect 50662 4678 50714 4730
rect 50714 4678 50716 4730
rect 50660 4676 50716 4678
rect 50764 4730 50820 4732
rect 50764 4678 50766 4730
rect 50766 4678 50818 4730
rect 50818 4678 50820 4730
rect 50764 4676 50820 4678
rect 8204 4508 8260 4564
rect 2492 3836 2548 3892
rect 4476 3946 4532 3948
rect 4476 3894 4478 3946
rect 4478 3894 4530 3946
rect 4530 3894 4532 3946
rect 4476 3892 4532 3894
rect 4580 3946 4636 3948
rect 4580 3894 4582 3946
rect 4582 3894 4634 3946
rect 4634 3894 4636 3946
rect 4580 3892 4636 3894
rect 4684 3946 4740 3948
rect 4684 3894 4686 3946
rect 4686 3894 4738 3946
rect 4738 3894 4740 3946
rect 4684 3892 4740 3894
rect 35196 3946 35252 3948
rect 35196 3894 35198 3946
rect 35198 3894 35250 3946
rect 35250 3894 35252 3946
rect 35196 3892 35252 3894
rect 35300 3946 35356 3948
rect 35300 3894 35302 3946
rect 35302 3894 35354 3946
rect 35354 3894 35356 3946
rect 35300 3892 35356 3894
rect 35404 3946 35460 3948
rect 35404 3894 35406 3946
rect 35406 3894 35458 3946
rect 35458 3894 35460 3946
rect 35404 3892 35460 3894
rect 1708 3276 1764 3332
rect 2716 3276 2772 3332
rect 19836 3162 19892 3164
rect 19836 3110 19838 3162
rect 19838 3110 19890 3162
rect 19890 3110 19892 3162
rect 19836 3108 19892 3110
rect 19940 3162 19996 3164
rect 19940 3110 19942 3162
rect 19942 3110 19994 3162
rect 19994 3110 19996 3162
rect 19940 3108 19996 3110
rect 20044 3162 20100 3164
rect 20044 3110 20046 3162
rect 20046 3110 20098 3162
rect 20098 3110 20100 3162
rect 20044 3108 20100 3110
rect 50556 3162 50612 3164
rect 50556 3110 50558 3162
rect 50558 3110 50610 3162
rect 50610 3110 50612 3162
rect 50556 3108 50612 3110
rect 50660 3162 50716 3164
rect 50660 3110 50662 3162
rect 50662 3110 50714 3162
rect 50714 3110 50716 3162
rect 50660 3108 50716 3110
rect 50764 3162 50820 3164
rect 50764 3110 50766 3162
rect 50766 3110 50818 3162
rect 50818 3110 50820 3162
rect 50764 3108 50820 3110
rect 1708 2044 1764 2100
<< metal3 >>
rect 0 57652 800 57680
rect 0 57596 2156 57652
rect 2212 57596 2222 57652
rect 0 57568 800 57596
rect 19826 56420 19836 56476
rect 19892 56420 19940 56476
rect 19996 56420 20044 56476
rect 20100 56420 20110 56476
rect 50546 56420 50556 56476
rect 50612 56420 50660 56476
rect 50716 56420 50764 56476
rect 50820 56420 50830 56476
rect 43250 56252 43260 56308
rect 43316 56252 44604 56308
rect 44660 56252 44670 56308
rect 47730 56252 47740 56308
rect 47796 56252 48972 56308
rect 49028 56252 49038 56308
rect 49970 56252 49980 56308
rect 50036 56252 52220 56308
rect 52276 56252 52286 56308
rect 54450 56252 54460 56308
rect 54516 56252 56028 56308
rect 56084 56252 56094 56308
rect 2146 56028 2156 56084
rect 2212 56028 2604 56084
rect 2660 56028 2670 56084
rect 27906 56028 27916 56084
rect 27972 56028 28588 56084
rect 28644 56028 28654 56084
rect 0 55860 800 55888
rect 0 55804 1708 55860
rect 1764 55804 3164 55860
rect 3220 55804 3230 55860
rect 30482 55804 30492 55860
rect 30548 55804 38892 55860
rect 38948 55804 40460 55860
rect 40516 55804 40526 55860
rect 0 55776 800 55804
rect 4466 55636 4476 55692
rect 4532 55636 4580 55692
rect 4636 55636 4684 55692
rect 4740 55636 4750 55692
rect 35186 55636 35196 55692
rect 35252 55636 35300 55692
rect 35356 55636 35404 55692
rect 35460 55636 35470 55692
rect 18498 55356 18508 55412
rect 18564 55356 20524 55412
rect 20580 55356 23212 55412
rect 23268 55356 23278 55412
rect 45490 55356 45500 55412
rect 45556 55356 46732 55412
rect 46788 55356 46798 55412
rect 52322 55356 52332 55412
rect 52388 55356 53676 55412
rect 53732 55356 53742 55412
rect 13570 55244 13580 55300
rect 13636 55244 16828 55300
rect 16884 55244 17724 55300
rect 17780 55244 21420 55300
rect 21476 55244 21486 55300
rect 29250 55244 29260 55300
rect 29316 55244 33180 55300
rect 33236 55244 33628 55300
rect 33684 55244 33694 55300
rect 5842 55132 5852 55188
rect 5908 55132 11788 55188
rect 11844 55132 11854 55188
rect 12674 55020 12684 55076
rect 12740 55020 15148 55076
rect 37090 55020 37100 55076
rect 37156 55020 37772 55076
rect 37828 55020 39900 55076
rect 39956 55020 40348 55076
rect 40404 55020 40414 55076
rect 15092 54740 15148 55020
rect 19826 54852 19836 54908
rect 19892 54852 19940 54908
rect 19996 54852 20044 54908
rect 20100 54852 20110 54908
rect 50546 54852 50556 54908
rect 50612 54852 50660 54908
rect 50716 54852 50764 54908
rect 50820 54852 50830 54908
rect 15092 54684 29148 54740
rect 29204 54684 29214 54740
rect 39106 54684 39116 54740
rect 39172 54684 40348 54740
rect 40404 54684 40796 54740
rect 40852 54684 41356 54740
rect 41412 54684 41422 54740
rect 1362 54572 1372 54628
rect 1428 54572 2044 54628
rect 2100 54572 2110 54628
rect 31826 54572 31836 54628
rect 31892 54572 36316 54628
rect 36372 54572 38220 54628
rect 38276 54572 38286 54628
rect 38882 54572 38892 54628
rect 38948 54572 41244 54628
rect 41300 54572 41692 54628
rect 41748 54572 41758 54628
rect 38220 54516 38276 54572
rect 17826 54460 17836 54516
rect 17892 54460 18396 54516
rect 18452 54460 18462 54516
rect 22866 54460 22876 54516
rect 22932 54460 23436 54516
rect 23492 54460 28812 54516
rect 28868 54460 30044 54516
rect 30100 54460 30110 54516
rect 38220 54460 40908 54516
rect 40964 54460 40974 54516
rect 24882 54348 24892 54404
rect 24948 54348 26012 54404
rect 26068 54348 26078 54404
rect 27570 54348 27580 54404
rect 27636 54348 32508 54404
rect 32564 54348 33404 54404
rect 33460 54348 33470 54404
rect 33954 54348 33964 54404
rect 34020 54348 36316 54404
rect 36372 54348 36382 54404
rect 29138 54236 29148 54292
rect 29204 54236 37884 54292
rect 37940 54236 37950 54292
rect 0 54068 800 54096
rect 4466 54068 4476 54124
rect 4532 54068 4580 54124
rect 4636 54068 4684 54124
rect 4740 54068 4750 54124
rect 35186 54068 35196 54124
rect 35252 54068 35300 54124
rect 35356 54068 35404 54124
rect 35460 54068 35470 54124
rect 0 54012 1708 54068
rect 1764 54012 2492 54068
rect 2548 54012 2558 54068
rect 0 53984 800 54012
rect 39442 53900 39452 53956
rect 39508 53900 43484 53956
rect 43540 53900 43550 53956
rect 2930 53788 2940 53844
rect 2996 53788 5740 53844
rect 5796 53788 5806 53844
rect 12786 53788 12796 53844
rect 12852 53788 16044 53844
rect 16100 53788 16110 53844
rect 22866 53788 22876 53844
rect 22932 53788 23660 53844
rect 23716 53788 23726 53844
rect 26562 53788 26572 53844
rect 26628 53788 28140 53844
rect 28196 53788 28206 53844
rect 30370 53788 30380 53844
rect 30436 53788 33292 53844
rect 33348 53788 33628 53844
rect 33684 53788 33694 53844
rect 39106 53788 39116 53844
rect 39172 53788 41692 53844
rect 41748 53788 41758 53844
rect 44594 53788 44604 53844
rect 44660 53788 54572 53844
rect 54628 53788 54638 53844
rect 21746 53676 21756 53732
rect 21812 53676 22428 53732
rect 22484 53676 22494 53732
rect 22642 53676 22652 53732
rect 22708 53676 27580 53732
rect 27636 53676 27646 53732
rect 32050 53676 32060 53732
rect 32116 53676 36988 53732
rect 37044 53676 37054 53732
rect 41234 53676 41244 53732
rect 41300 53676 43148 53732
rect 43204 53676 43214 53732
rect 22306 53564 22316 53620
rect 22372 53564 24556 53620
rect 24612 53564 24622 53620
rect 25218 53564 25228 53620
rect 25284 53564 26348 53620
rect 26404 53564 26414 53620
rect 31892 53564 32620 53620
rect 32676 53564 33068 53620
rect 33124 53564 34524 53620
rect 34580 53564 38444 53620
rect 38500 53564 38510 53620
rect 11554 53452 11564 53508
rect 11620 53452 18172 53508
rect 18228 53452 21980 53508
rect 22036 53452 22652 53508
rect 22708 53452 22718 53508
rect 24994 53452 25004 53508
rect 25060 53452 25676 53508
rect 25732 53452 29260 53508
rect 29316 53452 30268 53508
rect 30324 53452 30334 53508
rect 19826 53284 19836 53340
rect 19892 53284 19940 53340
rect 19996 53284 20044 53340
rect 20100 53284 20110 53340
rect 31892 53172 31948 53564
rect 50546 53284 50556 53340
rect 50612 53284 50660 53340
rect 50716 53284 50764 53340
rect 50820 53284 50830 53340
rect 12338 53116 12348 53172
rect 12404 53116 12796 53172
rect 12852 53116 13804 53172
rect 13860 53116 31948 53172
rect 34402 53116 34412 53172
rect 34468 53116 41020 53172
rect 41076 53116 41086 53172
rect 9874 53004 9884 53060
rect 9940 53004 10556 53060
rect 10612 53004 11116 53060
rect 11172 53004 11182 53060
rect 15474 53004 15484 53060
rect 15540 53004 22764 53060
rect 22820 53004 22830 53060
rect 23986 53004 23996 53060
rect 24052 53004 25452 53060
rect 25508 53004 26684 53060
rect 26740 53004 26750 53060
rect 30034 53004 30044 53060
rect 30100 53004 31948 53060
rect 32274 53004 32284 53060
rect 32340 53004 36764 53060
rect 36820 53004 36830 53060
rect 41570 53004 41580 53060
rect 41636 53004 41916 53060
rect 41972 53004 41982 53060
rect 31892 52948 31948 53004
rect 7970 52892 7980 52948
rect 8036 52892 10668 52948
rect 10724 52892 10734 52948
rect 10882 52892 10892 52948
rect 10948 52892 11564 52948
rect 11620 52892 11630 52948
rect 16146 52892 16156 52948
rect 16212 52892 17276 52948
rect 17332 52892 18060 52948
rect 18116 52892 18126 52948
rect 23538 52892 23548 52948
rect 23604 52892 26124 52948
rect 26180 52892 26190 52948
rect 31892 52892 33180 52948
rect 33236 52892 33246 52948
rect 33954 52892 33964 52948
rect 34020 52892 37772 52948
rect 37828 52892 37838 52948
rect 41458 52892 41468 52948
rect 41524 52892 42700 52948
rect 42756 52892 42766 52948
rect 1698 52780 1708 52836
rect 1764 52780 2492 52836
rect 2548 52780 2558 52836
rect 18162 52780 18172 52836
rect 18228 52780 19964 52836
rect 20020 52780 20030 52836
rect 21746 52780 21756 52836
rect 21812 52780 22540 52836
rect 22596 52780 22606 52836
rect 27010 52780 27020 52836
rect 27076 52780 27468 52836
rect 27524 52780 28476 52836
rect 28532 52780 28542 52836
rect 30818 52780 30828 52836
rect 30884 52780 31948 52836
rect 32004 52780 32014 52836
rect 36530 52780 36540 52836
rect 36596 52780 37660 52836
rect 37716 52780 37726 52836
rect 42578 52780 42588 52836
rect 42644 52780 44828 52836
rect 44884 52780 44894 52836
rect 27020 52724 27076 52780
rect 10434 52668 10444 52724
rect 10500 52668 11004 52724
rect 11060 52668 11676 52724
rect 11732 52668 11742 52724
rect 16482 52668 16492 52724
rect 16548 52668 27076 52724
rect 10210 52556 10220 52612
rect 10276 52556 12684 52612
rect 12740 52556 12750 52612
rect 15372 52556 24892 52612
rect 24948 52556 24958 52612
rect 4466 52500 4476 52556
rect 4532 52500 4580 52556
rect 4636 52500 4684 52556
rect 4740 52500 4750 52556
rect 15372 52500 15428 52556
rect 35186 52500 35196 52556
rect 35252 52500 35300 52556
rect 35356 52500 35404 52556
rect 35460 52500 35470 52556
rect 10322 52444 10332 52500
rect 10388 52444 12796 52500
rect 12852 52444 14812 52500
rect 14868 52444 15372 52500
rect 15428 52444 15438 52500
rect 17948 52444 18396 52500
rect 18452 52444 19068 52500
rect 19124 52444 25452 52500
rect 25508 52444 25518 52500
rect 17948 52388 18004 52444
rect 12348 52332 18004 52388
rect 0 52276 800 52304
rect 0 52220 1708 52276
rect 1764 52220 1774 52276
rect 0 52192 800 52220
rect 12348 52164 12404 52332
rect 14578 52220 14588 52276
rect 14644 52220 16156 52276
rect 16212 52220 16222 52276
rect 18050 52220 18060 52276
rect 18116 52220 19180 52276
rect 19236 52220 19246 52276
rect 23090 52220 23100 52276
rect 23156 52220 27244 52276
rect 27300 52220 27310 52276
rect 31892 52220 32844 52276
rect 32900 52220 32910 52276
rect 31892 52164 31948 52220
rect 11330 52108 11340 52164
rect 11396 52108 12348 52164
rect 12404 52108 12414 52164
rect 16258 52108 16268 52164
rect 16324 52108 16492 52164
rect 16548 52108 18620 52164
rect 18676 52108 18686 52164
rect 20626 52108 20636 52164
rect 20692 52108 21084 52164
rect 21140 52108 25228 52164
rect 25284 52108 29372 52164
rect 29428 52108 29438 52164
rect 29596 52108 31948 52164
rect 37426 52108 37436 52164
rect 37492 52108 38332 52164
rect 38388 52108 38398 52164
rect 29596 52052 29652 52108
rect 15586 51996 15596 52052
rect 15652 51996 17388 52052
rect 17444 51996 18172 52052
rect 18228 51996 18238 52052
rect 25442 51996 25452 52052
rect 25508 51996 26796 52052
rect 26852 51996 29596 52052
rect 29652 51996 29662 52052
rect 39218 51996 39228 52052
rect 39284 51996 42252 52052
rect 42308 51996 42318 52052
rect 3826 51884 3836 51940
rect 3892 51884 8428 51940
rect 8978 51884 8988 51940
rect 9044 51884 13244 51940
rect 13300 51884 13310 51940
rect 15138 51884 15148 51940
rect 15204 51884 15708 51940
rect 15764 51884 15774 51940
rect 8372 51828 8428 51884
rect 8372 51772 10108 51828
rect 10164 51772 10174 51828
rect 19826 51716 19836 51772
rect 19892 51716 19940 51772
rect 19996 51716 20044 51772
rect 20100 51716 20110 51772
rect 50546 51716 50556 51772
rect 50612 51716 50660 51772
rect 50716 51716 50764 51772
rect 50820 51716 50830 51772
rect 38098 51660 38108 51716
rect 38164 51660 40068 51716
rect 40012 51604 40068 51660
rect 10882 51548 10892 51604
rect 10948 51548 12012 51604
rect 12068 51548 15036 51604
rect 15092 51548 15102 51604
rect 17042 51548 17052 51604
rect 17108 51548 38668 51604
rect 38724 51548 38734 51604
rect 40002 51548 40012 51604
rect 40068 51548 42252 51604
rect 42308 51548 42318 51604
rect 2034 51436 2044 51492
rect 2100 51436 2716 51492
rect 2772 51436 2782 51492
rect 10770 51436 10780 51492
rect 10836 51436 11564 51492
rect 11620 51436 11630 51492
rect 37314 51436 37324 51492
rect 37380 51436 41244 51492
rect 41300 51436 41310 51492
rect 4386 51324 4396 51380
rect 4452 51324 5180 51380
rect 5236 51324 7644 51380
rect 7700 51324 8988 51380
rect 9044 51324 9054 51380
rect 26898 51324 26908 51380
rect 26964 51324 30492 51380
rect 30548 51324 30558 51380
rect 32498 51324 32508 51380
rect 32564 51324 38444 51380
rect 38500 51324 38510 51380
rect 38770 51324 38780 51380
rect 38836 51324 41020 51380
rect 41076 51324 41086 51380
rect 1810 51212 1820 51268
rect 1876 51212 2492 51268
rect 2548 51212 2558 51268
rect 5058 51212 5068 51268
rect 5124 51212 11900 51268
rect 11956 51212 11966 51268
rect 25890 51212 25900 51268
rect 25956 51212 27580 51268
rect 27636 51212 28252 51268
rect 28308 51212 28318 51268
rect 37874 51212 37884 51268
rect 37940 51212 38892 51268
rect 38948 51212 38958 51268
rect 15810 51100 15820 51156
rect 15876 51100 16828 51156
rect 16884 51100 17724 51156
rect 17780 51100 30380 51156
rect 30436 51100 30446 51156
rect 38434 51100 38444 51156
rect 38500 51100 39004 51156
rect 39060 51100 39070 51156
rect 39218 51100 39228 51156
rect 39284 51100 41580 51156
rect 41636 51100 41646 51156
rect 39004 51044 39060 51100
rect 39004 50988 40348 51044
rect 40404 50988 40414 51044
rect 4466 50932 4476 50988
rect 4532 50932 4580 50988
rect 4636 50932 4684 50988
rect 4740 50932 4750 50988
rect 35186 50932 35196 50988
rect 35252 50932 35300 50988
rect 35356 50932 35404 50988
rect 35460 50932 35470 50988
rect 5842 50764 5852 50820
rect 5908 50764 7308 50820
rect 7364 50764 7374 50820
rect 22418 50764 22428 50820
rect 22484 50764 26236 50820
rect 26292 50764 26302 50820
rect 26786 50764 26796 50820
rect 26852 50708 26908 50820
rect 1698 50652 1708 50708
rect 1764 50652 3276 50708
rect 3332 50652 3342 50708
rect 22978 50652 22988 50708
rect 23044 50652 23660 50708
rect 23716 50652 23726 50708
rect 26852 50652 27356 50708
rect 27412 50652 27422 50708
rect 37090 50652 37100 50708
rect 37156 50652 40460 50708
rect 40516 50652 40908 50708
rect 40964 50652 41244 50708
rect 41300 50652 41310 50708
rect 42466 50652 42476 50708
rect 42532 50652 44156 50708
rect 44212 50652 44222 50708
rect 15586 50540 15596 50596
rect 15652 50540 21868 50596
rect 21924 50540 24108 50596
rect 24164 50540 24444 50596
rect 24500 50540 24510 50596
rect 26002 50540 26012 50596
rect 26068 50540 26796 50596
rect 26852 50540 26862 50596
rect 0 50484 800 50512
rect 0 50428 1708 50484
rect 1764 50428 1774 50484
rect 13234 50428 13244 50484
rect 13300 50428 16492 50484
rect 16548 50428 17612 50484
rect 17668 50428 17678 50484
rect 23538 50428 23548 50484
rect 23604 50428 24556 50484
rect 24612 50428 24622 50484
rect 0 50400 800 50428
rect 17938 50316 17948 50372
rect 18004 50316 18284 50372
rect 18340 50316 18350 50372
rect 32386 50316 32396 50372
rect 32452 50316 32956 50372
rect 33012 50316 33516 50372
rect 33572 50316 37100 50372
rect 37156 50316 37166 50372
rect 19826 50148 19836 50204
rect 19892 50148 19940 50204
rect 19996 50148 20044 50204
rect 20100 50148 20110 50204
rect 50546 50148 50556 50204
rect 50612 50148 50660 50204
rect 50716 50148 50764 50204
rect 50820 50148 50830 50204
rect 11106 49980 11116 50036
rect 11172 49980 12012 50036
rect 12068 49980 12078 50036
rect 12562 49980 12572 50036
rect 12628 49980 13132 50036
rect 13188 49980 30380 50036
rect 30436 49980 30446 50036
rect 30706 49980 30716 50036
rect 30772 49980 33068 50036
rect 33124 49980 34076 50036
rect 34132 49980 34142 50036
rect 3826 49868 3836 49924
rect 3892 49868 10780 49924
rect 10836 49868 10846 49924
rect 17826 49868 17836 49924
rect 17892 49868 18396 49924
rect 18452 49868 22204 49924
rect 22260 49868 22270 49924
rect 23762 49868 23772 49924
rect 23828 49868 25228 49924
rect 25284 49868 25294 49924
rect 8978 49756 8988 49812
rect 9044 49756 10556 49812
rect 10612 49756 10622 49812
rect 29250 49756 29260 49812
rect 29316 49756 33292 49812
rect 33348 49756 33358 49812
rect 31826 49644 31836 49700
rect 31892 49644 33180 49700
rect 33236 49644 33246 49700
rect 34850 49644 34860 49700
rect 34916 49644 35644 49700
rect 35700 49644 35710 49700
rect 10546 49532 10556 49588
rect 10612 49532 11228 49588
rect 11284 49532 11294 49588
rect 33954 49532 33964 49588
rect 34020 49532 34300 49588
rect 34356 49532 34748 49588
rect 34804 49532 35420 49588
rect 35476 49532 35486 49588
rect 4466 49364 4476 49420
rect 4532 49364 4580 49420
rect 4636 49364 4684 49420
rect 4740 49364 4750 49420
rect 35186 49364 35196 49420
rect 35252 49364 35300 49420
rect 35356 49364 35404 49420
rect 35460 49364 35470 49420
rect 10098 49196 10108 49252
rect 10164 49196 11116 49252
rect 11172 49196 11182 49252
rect 26852 49084 29260 49140
rect 29316 49084 29326 49140
rect 8194 48972 8204 49028
rect 8260 48972 15372 49028
rect 15428 48972 15438 49028
rect 19058 48972 19068 49028
rect 19124 48972 21868 49028
rect 21924 48972 21934 49028
rect 24658 48972 24668 49028
rect 24724 48972 25564 49028
rect 25620 48972 25630 49028
rect 26852 48916 26908 49084
rect 7410 48860 7420 48916
rect 7476 48860 8092 48916
rect 8148 48860 8428 48916
rect 8484 48860 12796 48916
rect 12852 48860 12862 48916
rect 20402 48860 20412 48916
rect 20468 48860 26908 48916
rect 27122 48860 27132 48916
rect 27188 48860 45388 48916
rect 45444 48860 45454 48916
rect 10658 48748 10668 48804
rect 10724 48748 11340 48804
rect 11396 48748 11406 48804
rect 12450 48748 12460 48804
rect 12516 48748 12908 48804
rect 12964 48748 22036 48804
rect 36418 48748 36428 48804
rect 36484 48748 37156 48804
rect 0 48692 800 48720
rect 0 48636 1708 48692
rect 1764 48636 2492 48692
rect 2548 48636 2558 48692
rect 0 48608 800 48636
rect 19826 48580 19836 48636
rect 19892 48580 19940 48636
rect 19996 48580 20044 48636
rect 20100 48580 20110 48636
rect 8306 48412 8316 48468
rect 8372 48412 9660 48468
rect 9716 48412 9726 48468
rect 6626 48300 6636 48356
rect 6692 48300 7084 48356
rect 7140 48300 7150 48356
rect 10210 48300 10220 48356
rect 10276 48300 11452 48356
rect 11508 48300 11518 48356
rect 19590 48300 19628 48356
rect 19684 48300 19694 48356
rect 6066 48188 6076 48244
rect 6132 48188 10556 48244
rect 10612 48188 10622 48244
rect 16034 48188 16044 48244
rect 16100 48188 16492 48244
rect 16548 48188 20524 48244
rect 20580 48188 21644 48244
rect 21700 48188 21710 48244
rect 4466 47796 4476 47852
rect 4532 47796 4580 47852
rect 4636 47796 4684 47852
rect 4740 47796 4750 47852
rect 10556 47796 10612 48188
rect 21980 48132 22036 48748
rect 37100 48692 37156 48748
rect 22866 48636 22876 48692
rect 22932 48636 33516 48692
rect 33572 48636 34188 48692
rect 34244 48636 34254 48692
rect 37090 48636 37100 48692
rect 37156 48636 38556 48692
rect 38612 48636 40012 48692
rect 40068 48636 40078 48692
rect 50546 48580 50556 48636
rect 50612 48580 50660 48636
rect 50716 48580 50764 48636
rect 50820 48580 50830 48636
rect 31714 48524 31724 48580
rect 31780 48524 33068 48580
rect 33124 48524 33134 48580
rect 23202 48412 23212 48468
rect 23268 48412 23884 48468
rect 23940 48412 23950 48468
rect 22418 48300 22428 48356
rect 22484 48300 25788 48356
rect 25844 48300 25854 48356
rect 26002 48300 26012 48356
rect 26068 48300 29484 48356
rect 29540 48300 29550 48356
rect 31490 48300 31500 48356
rect 31556 48300 32172 48356
rect 32228 48300 32238 48356
rect 22194 48188 22204 48244
rect 22260 48188 22876 48244
rect 22932 48188 22942 48244
rect 23426 48188 23436 48244
rect 23492 48188 23996 48244
rect 24052 48188 24556 48244
rect 24612 48188 24622 48244
rect 26562 48188 26572 48244
rect 26628 48188 29036 48244
rect 29092 48188 29102 48244
rect 29810 48188 29820 48244
rect 29876 48188 39452 48244
rect 39508 48188 39518 48244
rect 14466 48076 14476 48132
rect 14532 48076 15260 48132
rect 15316 48076 15326 48132
rect 17602 48076 17612 48132
rect 17668 48076 18060 48132
rect 18116 48076 18620 48132
rect 18676 48076 19180 48132
rect 19236 48076 19246 48132
rect 21980 48076 26908 48132
rect 28578 48076 28588 48132
rect 28644 48076 32844 48132
rect 32900 48076 32910 48132
rect 11666 47964 11676 48020
rect 11732 47964 13916 48020
rect 13972 47964 13982 48020
rect 15810 47964 15820 48020
rect 15876 47964 22428 48020
rect 22484 47964 23436 48020
rect 23492 47964 23502 48020
rect 26852 47908 26908 48076
rect 29474 47964 29484 48020
rect 29540 47964 30940 48020
rect 30996 47964 31006 48020
rect 18274 47852 18284 47908
rect 18340 47852 18956 47908
rect 19012 47852 19022 47908
rect 21970 47852 21980 47908
rect 22036 47852 22540 47908
rect 22596 47852 22606 47908
rect 26852 47852 31500 47908
rect 31556 47852 31566 47908
rect 35186 47796 35196 47852
rect 35252 47796 35300 47852
rect 35356 47796 35404 47852
rect 35460 47796 35470 47852
rect 10556 47740 11340 47796
rect 11396 47740 11406 47796
rect 18610 47740 18620 47796
rect 18676 47740 23548 47796
rect 35746 47740 35756 47796
rect 35812 47740 37324 47796
rect 37380 47740 38332 47796
rect 38388 47740 38398 47796
rect 2146 47628 2156 47684
rect 2212 47628 3276 47684
rect 3332 47628 3342 47684
rect 13346 47628 13356 47684
rect 13412 47628 14476 47684
rect 14532 47628 14542 47684
rect 18498 47628 18508 47684
rect 18564 47628 18956 47684
rect 19012 47628 20076 47684
rect 20132 47628 20142 47684
rect 23492 47572 23548 47740
rect 24098 47628 24108 47684
rect 24164 47628 37772 47684
rect 37828 47628 37838 47684
rect 6402 47516 6412 47572
rect 6468 47516 11788 47572
rect 11844 47516 12124 47572
rect 12180 47516 12190 47572
rect 14242 47516 14252 47572
rect 14308 47516 16436 47572
rect 23492 47516 26908 47572
rect 32050 47516 32060 47572
rect 32116 47516 47740 47572
rect 47796 47516 47806 47572
rect 2482 47404 2492 47460
rect 2548 47404 3948 47460
rect 4004 47404 4014 47460
rect 8754 47404 8764 47460
rect 8820 47404 10780 47460
rect 10836 47404 10846 47460
rect 13122 47404 13132 47460
rect 13188 47404 14028 47460
rect 14084 47404 14812 47460
rect 14868 47404 14878 47460
rect 15362 47404 15372 47460
rect 15428 47404 16156 47460
rect 16212 47404 16222 47460
rect 15372 47348 15428 47404
rect 13570 47292 13580 47348
rect 13636 47292 14700 47348
rect 14756 47292 15428 47348
rect 16380 47348 16436 47516
rect 26852 47460 26908 47516
rect 17154 47404 17164 47460
rect 17220 47404 18284 47460
rect 18340 47404 20076 47460
rect 20132 47404 20142 47460
rect 26852 47404 27356 47460
rect 27412 47404 27422 47460
rect 27682 47404 27692 47460
rect 27748 47404 31276 47460
rect 31332 47404 31342 47460
rect 32834 47404 32844 47460
rect 32900 47404 33180 47460
rect 33236 47404 33246 47460
rect 34962 47404 34972 47460
rect 35028 47404 35756 47460
rect 35812 47404 35822 47460
rect 38098 47404 38108 47460
rect 38164 47404 38892 47460
rect 38948 47404 38958 47460
rect 40002 47404 40012 47460
rect 40068 47404 42700 47460
rect 42756 47404 42766 47460
rect 33180 47348 33236 47404
rect 16380 47292 31948 47348
rect 32004 47292 32014 47348
rect 33180 47292 38668 47348
rect 41234 47292 41244 47348
rect 41300 47292 42028 47348
rect 42084 47292 42094 47348
rect 38612 47236 38668 47292
rect 5730 47180 5740 47236
rect 5796 47180 24668 47236
rect 24724 47180 25228 47236
rect 25284 47180 25294 47236
rect 31154 47180 31164 47236
rect 31220 47180 33628 47236
rect 33684 47180 35084 47236
rect 35140 47180 35150 47236
rect 38612 47180 38780 47236
rect 38836 47180 38846 47236
rect 3714 47068 3724 47124
rect 3780 47068 4060 47124
rect 4116 47068 7308 47124
rect 7364 47068 8316 47124
rect 8372 47068 8382 47124
rect 14466 47068 14476 47124
rect 14532 47068 15484 47124
rect 15540 47068 16044 47124
rect 16100 47068 16110 47124
rect 18162 47068 18172 47124
rect 18228 47068 18620 47124
rect 18676 47068 18686 47124
rect 33282 47068 33292 47124
rect 33348 47068 33358 47124
rect 19826 47012 19836 47068
rect 19892 47012 19940 47068
rect 19996 47012 20044 47068
rect 20100 47012 20110 47068
rect 33292 47012 33348 47068
rect 50546 47012 50556 47068
rect 50612 47012 50660 47068
rect 50716 47012 50764 47068
rect 50820 47012 50830 47068
rect 22540 46956 26908 47012
rect 27906 46956 27916 47012
rect 27972 46956 33740 47012
rect 33796 46956 33806 47012
rect 38658 46956 38668 47012
rect 38724 46956 39228 47012
rect 39284 46956 39788 47012
rect 39844 46956 39854 47012
rect 40338 46956 40348 47012
rect 40404 46956 41132 47012
rect 41188 46956 41198 47012
rect 0 46900 800 46928
rect 22540 46900 22596 46956
rect 26852 46900 26908 46956
rect 0 46844 1708 46900
rect 1764 46844 2492 46900
rect 2548 46844 2558 46900
rect 4498 46844 4508 46900
rect 4564 46844 8988 46900
rect 9044 46844 10332 46900
rect 10388 46844 10398 46900
rect 12898 46844 12908 46900
rect 12964 46844 13356 46900
rect 13412 46844 13422 46900
rect 22530 46844 22540 46900
rect 22596 46844 22606 46900
rect 23986 46844 23996 46900
rect 24052 46844 24892 46900
rect 24948 46844 24958 46900
rect 26852 46844 29596 46900
rect 29652 46844 29662 46900
rect 32722 46844 32732 46900
rect 32788 46844 34076 46900
rect 34132 46844 34860 46900
rect 34916 46844 34926 46900
rect 39106 46844 39116 46900
rect 39172 46844 40908 46900
rect 40964 46844 40974 46900
rect 0 46816 800 46844
rect 4834 46732 4844 46788
rect 4900 46732 7868 46788
rect 7924 46732 9100 46788
rect 9156 46732 9166 46788
rect 12786 46732 12796 46788
rect 12852 46732 13132 46788
rect 13188 46732 13198 46788
rect 13804 46732 28812 46788
rect 28868 46732 28878 46788
rect 35186 46732 35196 46788
rect 35252 46732 36652 46788
rect 36708 46732 36718 46788
rect 38434 46732 38444 46788
rect 38500 46732 39564 46788
rect 39620 46732 41468 46788
rect 41524 46732 41534 46788
rect 7522 46620 7532 46676
rect 7588 46620 7756 46676
rect 7812 46620 11452 46676
rect 11508 46620 11518 46676
rect 13804 46564 13860 46732
rect 14018 46620 14028 46676
rect 14084 46620 15036 46676
rect 15092 46620 15102 46676
rect 20066 46620 20076 46676
rect 20132 46620 21308 46676
rect 21364 46620 21374 46676
rect 26852 46620 31164 46676
rect 31220 46620 31230 46676
rect 32610 46620 32620 46676
rect 32676 46620 33292 46676
rect 33348 46620 33358 46676
rect 12562 46508 12572 46564
rect 12628 46508 13860 46564
rect 15036 46564 15092 46620
rect 15036 46508 15148 46564
rect 19618 46508 19628 46564
rect 19684 46508 21756 46564
rect 21812 46508 21822 46564
rect 15092 46452 15148 46508
rect 26852 46452 26908 46620
rect 30370 46508 30380 46564
rect 30436 46508 32508 46564
rect 32564 46508 32574 46564
rect 15092 46396 15708 46452
rect 15764 46396 16380 46452
rect 16436 46396 26908 46452
rect 29586 46396 29596 46452
rect 29652 46396 32956 46452
rect 33012 46396 33022 46452
rect 20972 46284 29260 46340
rect 29316 46284 29326 46340
rect 4466 46228 4476 46284
rect 4532 46228 4580 46284
rect 4636 46228 4684 46284
rect 4740 46228 4750 46284
rect 14466 46060 14476 46116
rect 14532 46060 15820 46116
rect 15876 46060 15886 46116
rect 20972 46004 21028 46284
rect 35186 46228 35196 46284
rect 35252 46228 35300 46284
rect 35356 46228 35404 46284
rect 35460 46228 35470 46284
rect 22642 46172 22652 46228
rect 22708 46172 34524 46228
rect 34580 46172 34590 46228
rect 23622 46060 23660 46116
rect 23716 46060 23726 46116
rect 28242 46060 28252 46116
rect 28308 46060 29372 46116
rect 29428 46060 29438 46116
rect 9874 45948 9884 46004
rect 9940 45948 11004 46004
rect 11060 45948 12012 46004
rect 12068 45948 12078 46004
rect 15092 45948 21028 46004
rect 32050 45948 32060 46004
rect 32116 45948 50316 46004
rect 50372 45948 50382 46004
rect 15092 45892 15148 45948
rect 8642 45836 8652 45892
rect 8708 45836 9548 45892
rect 9604 45836 10892 45892
rect 10948 45836 10958 45892
rect 11116 45836 15148 45892
rect 16706 45836 16716 45892
rect 16772 45836 17388 45892
rect 17444 45836 17454 45892
rect 20290 45836 20300 45892
rect 20356 45836 21420 45892
rect 21476 45836 21486 45892
rect 26758 45836 26796 45892
rect 26852 45836 26862 45892
rect 31826 45836 31836 45892
rect 31892 45836 38556 45892
rect 38612 45836 38622 45892
rect 11116 45780 11172 45836
rect 4498 45724 4508 45780
rect 4564 45724 8764 45780
rect 8820 45724 9324 45780
rect 9380 45724 9390 45780
rect 9548 45724 11172 45780
rect 11330 45724 11340 45780
rect 11396 45724 12124 45780
rect 12180 45724 12190 45780
rect 16482 45724 16492 45780
rect 16548 45724 17836 45780
rect 17892 45724 21084 45780
rect 21140 45724 21150 45780
rect 24546 45724 24556 45780
rect 24612 45724 27356 45780
rect 27412 45724 27422 45780
rect 33506 45724 33516 45780
rect 33572 45724 34188 45780
rect 34244 45724 34254 45780
rect 40226 45724 40236 45780
rect 40292 45724 41356 45780
rect 41412 45724 41422 45780
rect 9548 45668 9604 45724
rect 7074 45612 7084 45668
rect 7140 45612 8092 45668
rect 8148 45612 8158 45668
rect 8306 45612 8316 45668
rect 8372 45612 9604 45668
rect 10434 45612 10444 45668
rect 10500 45612 10556 45668
rect 10612 45612 10622 45668
rect 10770 45612 10780 45668
rect 10836 45612 11452 45668
rect 11508 45612 11518 45668
rect 15092 45612 28364 45668
rect 28420 45612 28430 45668
rect 33394 45612 33404 45668
rect 33460 45612 34524 45668
rect 34580 45612 34590 45668
rect 6178 45500 6188 45556
rect 6244 45500 6972 45556
rect 7028 45500 7038 45556
rect 15092 45444 15148 45612
rect 18834 45500 18844 45556
rect 18900 45500 19628 45556
rect 19684 45500 19694 45556
rect 20178 45500 20188 45556
rect 20244 45500 21420 45556
rect 21476 45500 22764 45556
rect 22820 45500 22830 45556
rect 27122 45500 27132 45556
rect 27188 45500 28140 45556
rect 28196 45500 28206 45556
rect 4162 45388 4172 45444
rect 4228 45388 6524 45444
rect 6580 45388 6748 45444
rect 6804 45388 7980 45444
rect 8036 45388 8046 45444
rect 8204 45388 15148 45444
rect 8204 45332 8260 45388
rect 4050 45276 4060 45332
rect 4116 45276 8260 45332
rect 19628 45332 19684 45500
rect 19826 45444 19836 45500
rect 19892 45444 19940 45500
rect 19996 45444 20044 45500
rect 20100 45444 20110 45500
rect 50546 45444 50556 45500
rect 50612 45444 50660 45500
rect 50716 45444 50764 45500
rect 50820 45444 50830 45500
rect 21186 45388 21196 45444
rect 21252 45388 23100 45444
rect 23156 45388 23166 45444
rect 19628 45276 20748 45332
rect 20804 45276 20814 45332
rect 23426 45276 23436 45332
rect 23492 45276 29372 45332
rect 29428 45276 29438 45332
rect 23650 45164 23660 45220
rect 23716 45164 24668 45220
rect 24724 45164 24734 45220
rect 25890 45164 25900 45220
rect 25956 45164 28700 45220
rect 28756 45164 28766 45220
rect 0 45108 800 45136
rect 0 45052 1708 45108
rect 1764 45052 2268 45108
rect 2324 45052 2334 45108
rect 2482 45052 2492 45108
rect 2548 45052 3052 45108
rect 3108 45052 3118 45108
rect 7746 45052 7756 45108
rect 7812 45052 13804 45108
rect 13860 45052 13870 45108
rect 17714 45052 17724 45108
rect 17780 45052 26124 45108
rect 26180 45052 26190 45108
rect 39442 45052 39452 45108
rect 39508 45052 40348 45108
rect 40404 45052 40414 45108
rect 0 45024 800 45052
rect 16258 44940 16268 44996
rect 16324 44940 20300 44996
rect 20356 44940 20860 44996
rect 20916 44940 20926 44996
rect 24322 44940 24332 44996
rect 24388 44940 25564 44996
rect 25620 44940 25630 44996
rect 37538 44940 37548 44996
rect 37604 44940 40124 44996
rect 40180 44940 44492 44996
rect 44548 44940 44558 44996
rect 1474 44828 1484 44884
rect 1540 44828 3164 44884
rect 3220 44828 3230 44884
rect 10434 44828 10444 44884
rect 10500 44828 11228 44884
rect 11284 44828 11294 44884
rect 17378 44828 17388 44884
rect 17444 44828 19292 44884
rect 19348 44828 19358 44884
rect 10546 44716 10556 44772
rect 10612 44716 11116 44772
rect 11172 44716 11182 44772
rect 4466 44660 4476 44716
rect 4532 44660 4580 44716
rect 4636 44660 4684 44716
rect 4740 44660 4750 44716
rect 35186 44660 35196 44716
rect 35252 44660 35300 44716
rect 35356 44660 35404 44716
rect 35460 44660 35470 44716
rect 14802 44604 14812 44660
rect 14868 44604 18844 44660
rect 18900 44604 18910 44660
rect 19954 44604 19964 44660
rect 20020 44604 21644 44660
rect 21700 44604 22988 44660
rect 23044 44604 23212 44660
rect 23268 44604 23278 44660
rect 24322 44604 24332 44660
rect 24388 44604 24668 44660
rect 24724 44604 26348 44660
rect 26404 44604 26414 44660
rect 14466 44492 14476 44548
rect 14532 44492 18620 44548
rect 18676 44492 20972 44548
rect 21028 44492 21038 44548
rect 21746 44492 21756 44548
rect 21812 44492 22092 44548
rect 22148 44492 22158 44548
rect 24668 44492 30156 44548
rect 30212 44492 30222 44548
rect 32162 44492 32172 44548
rect 32228 44492 34748 44548
rect 34804 44492 35420 44548
rect 35476 44492 40796 44548
rect 40852 44492 40862 44548
rect 24668 44436 24724 44492
rect 13010 44380 13020 44436
rect 13076 44380 15148 44436
rect 17490 44380 17500 44436
rect 17556 44380 19628 44436
rect 19684 44380 20524 44436
rect 20580 44380 20590 44436
rect 24658 44380 24668 44436
rect 24724 44380 24734 44436
rect 26114 44380 26124 44436
rect 26180 44380 26236 44436
rect 26292 44380 27020 44436
rect 27076 44380 27086 44436
rect 32722 44380 32732 44436
rect 32788 44380 55356 44436
rect 55412 44380 55422 44436
rect 15092 44324 15148 44380
rect 7970 44268 7980 44324
rect 8036 44268 10444 44324
rect 10500 44268 11004 44324
rect 11060 44268 11070 44324
rect 15092 44268 16604 44324
rect 16660 44268 16670 44324
rect 16818 44268 16828 44324
rect 16884 44268 18060 44324
rect 18116 44268 18126 44324
rect 20738 44268 20748 44324
rect 20804 44268 23436 44324
rect 23492 44268 23502 44324
rect 24546 44268 24556 44324
rect 24612 44268 26684 44324
rect 26740 44268 26750 44324
rect 30034 44268 30044 44324
rect 30100 44268 30828 44324
rect 30884 44268 30894 44324
rect 33506 44268 33516 44324
rect 33572 44268 34188 44324
rect 34244 44268 34254 44324
rect 36306 44268 36316 44324
rect 36372 44268 38556 44324
rect 38612 44268 39116 44324
rect 39172 44268 39182 44324
rect 6850 44156 6860 44212
rect 6916 44156 8092 44212
rect 8148 44156 8158 44212
rect 16930 44156 16940 44212
rect 16996 44156 17388 44212
rect 17444 44156 17454 44212
rect 18722 44156 18732 44212
rect 18788 44156 19852 44212
rect 19908 44156 21868 44212
rect 21924 44156 21934 44212
rect 22642 44156 22652 44212
rect 22708 44156 23660 44212
rect 23716 44156 24220 44212
rect 24276 44156 26460 44212
rect 26516 44156 26526 44212
rect 28466 44156 28476 44212
rect 28532 44156 31724 44212
rect 31780 44156 32956 44212
rect 33012 44156 33022 44212
rect 33282 44156 33292 44212
rect 33348 44156 37436 44212
rect 37492 44156 37502 44212
rect 2258 44044 2268 44100
rect 2324 44044 2716 44100
rect 2772 44044 2782 44100
rect 17266 44044 17276 44100
rect 17332 44044 17724 44100
rect 17780 44044 17790 44100
rect 19282 44044 19292 44100
rect 19348 44044 23100 44100
rect 23156 44044 23166 44100
rect 24994 44044 25004 44100
rect 25060 44044 27468 44100
rect 27524 44044 27534 44100
rect 9986 43932 9996 43988
rect 10052 43932 12684 43988
rect 12740 43932 12750 43988
rect 15698 43932 15708 43988
rect 15764 43932 16268 43988
rect 16324 43932 16334 43988
rect 26338 43932 26348 43988
rect 26404 43932 29148 43988
rect 29204 43932 29214 43988
rect 19826 43876 19836 43932
rect 19892 43876 19940 43932
rect 19996 43876 20044 43932
rect 20100 43876 20110 43932
rect 50546 43876 50556 43932
rect 50612 43876 50660 43932
rect 50716 43876 50764 43932
rect 50820 43876 50830 43932
rect 10546 43820 10556 43876
rect 10612 43820 19684 43876
rect 23762 43820 23772 43876
rect 23828 43820 24556 43876
rect 24612 43820 24622 43876
rect 6850 43708 6860 43764
rect 6916 43708 7308 43764
rect 7364 43708 7980 43764
rect 8036 43708 8046 43764
rect 8530 43708 8540 43764
rect 8596 43708 11340 43764
rect 11396 43708 11676 43764
rect 11732 43708 11742 43764
rect 12674 43708 12684 43764
rect 12740 43708 15260 43764
rect 15316 43708 15596 43764
rect 15652 43708 15662 43764
rect 16370 43708 16380 43764
rect 16436 43708 17500 43764
rect 17556 43708 17566 43764
rect 19628 43652 19684 43820
rect 22306 43708 22316 43764
rect 22372 43708 30604 43764
rect 30660 43708 30670 43764
rect 2034 43596 2044 43652
rect 2100 43596 2110 43652
rect 2706 43596 2716 43652
rect 2772 43596 2782 43652
rect 3602 43596 3612 43652
rect 3668 43596 4844 43652
rect 4900 43596 5292 43652
rect 5348 43596 6524 43652
rect 6580 43596 6590 43652
rect 7746 43596 7756 43652
rect 7812 43596 11004 43652
rect 11060 43596 12124 43652
rect 12180 43596 13132 43652
rect 13188 43596 13198 43652
rect 17602 43596 17612 43652
rect 17668 43596 19068 43652
rect 19124 43596 19134 43652
rect 19628 43596 23548 43652
rect 23604 43596 23614 43652
rect 23986 43596 23996 43652
rect 24052 43596 26572 43652
rect 26628 43596 26638 43652
rect 26852 43596 29148 43652
rect 29204 43596 29214 43652
rect 31714 43596 31724 43652
rect 31780 43596 32620 43652
rect 32676 43596 33068 43652
rect 33124 43596 33134 43652
rect 33394 43596 33404 43652
rect 33460 43596 34972 43652
rect 35028 43596 35038 43652
rect 39442 43596 39452 43652
rect 39508 43596 39676 43652
rect 39732 43596 41692 43652
rect 41748 43596 41758 43652
rect 2044 43540 2100 43596
rect 2044 43484 2380 43540
rect 2436 43484 2446 43540
rect 2716 43428 2772 43596
rect 26852 43540 26908 43596
rect 10098 43484 10108 43540
rect 10164 43484 13916 43540
rect 13972 43484 13982 43540
rect 16594 43484 16604 43540
rect 16660 43484 18620 43540
rect 18676 43484 18686 43540
rect 24210 43484 24220 43540
rect 24276 43484 26908 43540
rect 36978 43484 36988 43540
rect 37044 43484 40012 43540
rect 40068 43484 41020 43540
rect 41076 43484 41580 43540
rect 41636 43484 41646 43540
rect 2034 43372 2044 43428
rect 2100 43372 2772 43428
rect 4050 43372 4060 43428
rect 4116 43372 7868 43428
rect 7924 43372 7934 43428
rect 9986 43372 9996 43428
rect 10052 43372 11788 43428
rect 11844 43372 11854 43428
rect 12114 43372 12124 43428
rect 12180 43372 12460 43428
rect 12516 43372 12526 43428
rect 0 43316 800 43344
rect 13468 43316 13524 43484
rect 23062 43372 23100 43428
rect 23156 43372 25564 43428
rect 25620 43372 25630 43428
rect 29922 43372 29932 43428
rect 29988 43372 31052 43428
rect 31108 43372 31118 43428
rect 37202 43372 37212 43428
rect 37268 43372 38668 43428
rect 38724 43372 38734 43428
rect 40226 43372 40236 43428
rect 40292 43372 41132 43428
rect 41188 43372 41198 43428
rect 0 43260 1820 43316
rect 1876 43260 1886 43316
rect 3714 43260 3724 43316
rect 3780 43260 4508 43316
rect 4564 43260 11452 43316
rect 11508 43260 11900 43316
rect 11956 43260 11966 43316
rect 13458 43260 13468 43316
rect 13524 43260 13534 43316
rect 21746 43260 21756 43316
rect 21812 43260 24220 43316
rect 24276 43260 24286 43316
rect 24658 43260 24668 43316
rect 24724 43260 24734 43316
rect 33506 43260 33516 43316
rect 33572 43260 36428 43316
rect 36484 43260 36494 43316
rect 0 43232 800 43260
rect 24668 43204 24724 43260
rect 24668 43148 28588 43204
rect 28644 43148 28654 43204
rect 4466 43092 4476 43148
rect 4532 43092 4580 43148
rect 4636 43092 4684 43148
rect 4740 43092 4750 43148
rect 35186 43092 35196 43148
rect 35252 43092 35300 43148
rect 35356 43092 35404 43148
rect 35460 43092 35470 43148
rect 10434 43036 10444 43092
rect 10500 43036 11340 43092
rect 11396 43036 11406 43092
rect 12674 43036 12684 43092
rect 12740 43036 24108 43092
rect 24164 43036 24174 43092
rect 3332 42924 18732 42980
rect 18788 42924 18798 42980
rect 34402 42924 34412 42980
rect 34468 42924 35308 42980
rect 35364 42924 35374 42980
rect 3332 42532 3388 42924
rect 8306 42812 8316 42868
rect 8372 42812 21084 42868
rect 21140 42812 21150 42868
rect 23202 42812 23212 42868
rect 23268 42812 23884 42868
rect 23940 42812 23950 42868
rect 38658 42812 38668 42868
rect 38724 42812 39228 42868
rect 39284 42812 39294 42868
rect 41346 42812 41356 42868
rect 41412 42812 44044 42868
rect 44100 42812 44110 42868
rect 7858 42700 7868 42756
rect 7924 42700 8764 42756
rect 8820 42700 9324 42756
rect 9380 42700 9390 42756
rect 9762 42700 9772 42756
rect 9828 42700 10780 42756
rect 10836 42700 10846 42756
rect 16706 42700 16716 42756
rect 16772 42700 17052 42756
rect 17108 42700 17612 42756
rect 17668 42700 17678 42756
rect 18508 42700 24444 42756
rect 24500 42700 25004 42756
rect 25060 42700 25564 42756
rect 25620 42700 25630 42756
rect 28242 42700 28252 42756
rect 28308 42700 29372 42756
rect 29428 42700 29438 42756
rect 33506 42700 33516 42756
rect 33572 42700 38556 42756
rect 38612 42700 38622 42756
rect 18508 42644 18564 42700
rect 8194 42588 8204 42644
rect 8260 42588 8876 42644
rect 8932 42588 8942 42644
rect 10882 42588 10892 42644
rect 10948 42588 11788 42644
rect 11844 42588 11854 42644
rect 15138 42588 15148 42644
rect 15204 42588 18564 42644
rect 18722 42588 18732 42644
rect 18788 42588 25452 42644
rect 25508 42588 27916 42644
rect 27972 42588 27982 42644
rect 38994 42588 39004 42644
rect 39060 42588 40236 42644
rect 40292 42588 40302 42644
rect 40450 42588 40460 42644
rect 40516 42588 41916 42644
rect 41972 42588 41982 42644
rect 3042 42476 3052 42532
rect 3108 42476 3388 42532
rect 10210 42476 10220 42532
rect 10276 42476 10332 42532
rect 10388 42476 10398 42532
rect 18050 42476 18060 42532
rect 18116 42476 21308 42532
rect 21364 42476 21374 42532
rect 23090 42476 23100 42532
rect 23156 42476 23660 42532
rect 23716 42476 23996 42532
rect 24052 42476 24062 42532
rect 26786 42476 26796 42532
rect 26852 42476 30268 42532
rect 30324 42476 30334 42532
rect 32834 42476 32844 42532
rect 32900 42476 38668 42532
rect 38612 42420 38668 42476
rect 11330 42364 11340 42420
rect 11396 42364 17836 42420
rect 17892 42364 17902 42420
rect 20738 42364 20748 42420
rect 20804 42364 21868 42420
rect 21924 42364 21934 42420
rect 23846 42364 23884 42420
rect 23940 42364 23950 42420
rect 24658 42364 24668 42420
rect 24724 42364 25452 42420
rect 25508 42364 25518 42420
rect 33954 42364 33964 42420
rect 34020 42364 36988 42420
rect 37044 42364 37054 42420
rect 38612 42364 44604 42420
rect 44660 42364 44670 42420
rect 19826 42308 19836 42364
rect 19892 42308 19940 42364
rect 19996 42308 20044 42364
rect 20100 42308 20110 42364
rect 50546 42308 50556 42364
rect 50612 42308 50660 42364
rect 50716 42308 50764 42364
rect 50820 42308 50830 42364
rect 2706 42252 2716 42308
rect 2772 42252 3052 42308
rect 3108 42252 3118 42308
rect 5842 42252 5852 42308
rect 5908 42252 6636 42308
rect 6692 42252 9660 42308
rect 9716 42252 9726 42308
rect 12226 42252 12236 42308
rect 12292 42252 13804 42308
rect 13860 42252 13870 42308
rect 23650 42252 23660 42308
rect 23716 42252 24220 42308
rect 24276 42252 24286 42308
rect 8866 42140 8876 42196
rect 8932 42140 14252 42196
rect 14308 42140 15148 42196
rect 22866 42140 22876 42196
rect 22932 42140 30828 42196
rect 30884 42140 30894 42196
rect 15092 42084 15148 42140
rect 6402 42028 6412 42084
rect 6468 42028 7196 42084
rect 7252 42028 7644 42084
rect 7700 42028 7710 42084
rect 15092 42028 18060 42084
rect 18116 42028 18126 42084
rect 27346 42028 27356 42084
rect 27412 42028 32844 42084
rect 32900 42028 32910 42084
rect 34626 42028 34636 42084
rect 34692 42028 35196 42084
rect 35252 42028 35262 42084
rect 2034 41916 2044 41972
rect 2100 41916 2716 41972
rect 2772 41916 2782 41972
rect 16594 41916 16604 41972
rect 16660 41916 17948 41972
rect 18004 41916 18014 41972
rect 18162 41916 18172 41972
rect 18228 41916 20188 41972
rect 20244 41916 20254 41972
rect 20962 41916 20972 41972
rect 21028 41916 21980 41972
rect 22036 41916 22046 41972
rect 29586 41916 29596 41972
rect 29652 41916 30156 41972
rect 30212 41916 30222 41972
rect 32050 41916 32060 41972
rect 32116 41916 33516 41972
rect 33572 41916 34524 41972
rect 34580 41916 34590 41972
rect 35410 41916 35420 41972
rect 35476 41916 37772 41972
rect 37828 41916 37838 41972
rect 4050 41804 4060 41860
rect 4116 41804 6748 41860
rect 6804 41804 6814 41860
rect 9426 41804 9436 41860
rect 9492 41804 21532 41860
rect 21588 41804 22204 41860
rect 22260 41804 22270 41860
rect 23314 41804 23324 41860
rect 23380 41804 26572 41860
rect 26628 41804 26908 41860
rect 26964 41804 26974 41860
rect 34066 41804 34076 41860
rect 34132 41804 35084 41860
rect 35140 41804 39900 41860
rect 39956 41804 40460 41860
rect 40516 41804 40526 41860
rect 18834 41692 18844 41748
rect 18900 41692 19516 41748
rect 19572 41692 19582 41748
rect 21970 41692 21980 41748
rect 22036 41692 23436 41748
rect 23492 41692 23502 41748
rect 25330 41692 25340 41748
rect 25396 41692 27132 41748
rect 27188 41692 27804 41748
rect 27860 41692 28364 41748
rect 28420 41692 28430 41748
rect 34626 41692 34636 41748
rect 34692 41692 35756 41748
rect 35812 41692 35822 41748
rect 19282 41580 19292 41636
rect 19348 41580 19852 41636
rect 19908 41580 20636 41636
rect 20692 41580 20702 41636
rect 20850 41580 20860 41636
rect 20916 41580 23212 41636
rect 23268 41580 23278 41636
rect 0 41524 800 41552
rect 4466 41524 4476 41580
rect 4532 41524 4580 41580
rect 4636 41524 4684 41580
rect 4740 41524 4750 41580
rect 35186 41524 35196 41580
rect 35252 41524 35300 41580
rect 35356 41524 35404 41580
rect 35460 41524 35470 41580
rect 0 41468 1708 41524
rect 1764 41468 1774 41524
rect 21970 41468 21980 41524
rect 22036 41468 24668 41524
rect 24724 41468 24734 41524
rect 0 41440 800 41468
rect 14914 41356 14924 41412
rect 14980 41356 20188 41412
rect 20244 41356 20254 41412
rect 20850 41356 20860 41412
rect 20916 41356 21756 41412
rect 21812 41356 21822 41412
rect 23090 41356 23100 41412
rect 23156 41356 24892 41412
rect 24948 41356 24958 41412
rect 35298 41356 35308 41412
rect 35364 41356 35644 41412
rect 35700 41356 35710 41412
rect 9538 41244 9548 41300
rect 9604 41244 9884 41300
rect 9940 41244 9950 41300
rect 13010 41244 13020 41300
rect 13076 41244 27916 41300
rect 27972 41244 27982 41300
rect 2594 41132 2604 41188
rect 2660 41132 4060 41188
rect 4116 41132 4126 41188
rect 14018 41132 14028 41188
rect 14084 41132 15036 41188
rect 15092 41132 15102 41188
rect 15484 41132 16212 41188
rect 16370 41132 16380 41188
rect 16436 41132 17612 41188
rect 17668 41132 17678 41188
rect 19506 41132 19516 41188
rect 19572 41132 20804 41188
rect 21410 41132 21420 41188
rect 21476 41132 21756 41188
rect 21812 41132 21822 41188
rect 22204 41132 27020 41188
rect 27076 41132 27086 41188
rect 28466 41132 28476 41188
rect 28532 41132 29596 41188
rect 29652 41132 29662 41188
rect 33506 41132 33516 41188
rect 33572 41132 40908 41188
rect 40964 41132 40974 41188
rect 15484 41076 15540 41132
rect 2482 41020 2492 41076
rect 2548 41020 2716 41076
rect 2772 41020 2782 41076
rect 9538 41020 9548 41076
rect 9604 41020 13580 41076
rect 13636 41020 13646 41076
rect 14130 41020 14140 41076
rect 14196 41020 15540 41076
rect 16156 41076 16212 41132
rect 20748 41076 20804 41132
rect 22204 41076 22260 41132
rect 16156 41020 19852 41076
rect 19908 41020 20524 41076
rect 20580 41020 20590 41076
rect 20748 41020 22260 41076
rect 22530 41020 22540 41076
rect 22596 41020 23324 41076
rect 23380 41020 23390 41076
rect 26450 41020 26460 41076
rect 26516 41020 31052 41076
rect 31108 41020 31118 41076
rect 12226 40908 12236 40964
rect 12292 40908 27356 40964
rect 27412 40908 27422 40964
rect 29138 40908 29148 40964
rect 29204 40908 30380 40964
rect 30436 40908 30446 40964
rect 33058 40908 33068 40964
rect 33124 40908 52108 40964
rect 52164 40908 52174 40964
rect 12114 40796 12124 40852
rect 12180 40796 15708 40852
rect 15764 40796 15774 40852
rect 27122 40796 27132 40852
rect 27188 40796 27692 40852
rect 27748 40796 30044 40852
rect 30100 40796 30110 40852
rect 19826 40740 19836 40796
rect 19892 40740 19940 40796
rect 19996 40740 20044 40796
rect 20100 40740 20110 40796
rect 50546 40740 50556 40796
rect 50612 40740 50660 40796
rect 50716 40740 50764 40796
rect 50820 40740 50830 40796
rect 10546 40684 10556 40740
rect 10612 40684 11452 40740
rect 11508 40684 11518 40740
rect 13346 40684 13356 40740
rect 13412 40684 16156 40740
rect 16212 40684 16222 40740
rect 17490 40684 17500 40740
rect 17556 40684 18284 40740
rect 18340 40684 18350 40740
rect 27570 40684 27580 40740
rect 27636 40684 28588 40740
rect 28644 40684 28654 40740
rect 34066 40684 34076 40740
rect 34132 40684 34524 40740
rect 34580 40684 36092 40740
rect 36148 40684 36158 40740
rect 6626 40572 6636 40628
rect 6692 40572 18172 40628
rect 18228 40572 18732 40628
rect 18788 40572 18798 40628
rect 20178 40572 20188 40628
rect 20244 40572 21084 40628
rect 21140 40572 21980 40628
rect 22036 40572 22046 40628
rect 23202 40572 23212 40628
rect 23268 40572 25116 40628
rect 25172 40572 25182 40628
rect 27346 40572 27356 40628
rect 27412 40572 29484 40628
rect 29540 40572 29550 40628
rect 34626 40572 34636 40628
rect 34692 40572 35308 40628
rect 35364 40572 35374 40628
rect 4946 40460 4956 40516
rect 5012 40460 6188 40516
rect 6244 40460 6254 40516
rect 7186 40460 7196 40516
rect 7252 40460 8764 40516
rect 8820 40460 8830 40516
rect 9874 40460 9884 40516
rect 9940 40460 11676 40516
rect 11732 40460 11742 40516
rect 15250 40460 15260 40516
rect 15316 40460 17500 40516
rect 17556 40460 17566 40516
rect 18946 40460 18956 40516
rect 19012 40460 22316 40516
rect 22372 40460 22382 40516
rect 22540 40460 23884 40516
rect 23940 40460 23950 40516
rect 26114 40460 26124 40516
rect 26180 40460 26348 40516
rect 26404 40460 27244 40516
rect 27300 40460 27310 40516
rect 27794 40460 27804 40516
rect 27860 40460 31276 40516
rect 31332 40460 31342 40516
rect 22540 40404 22596 40460
rect 5058 40348 5068 40404
rect 5124 40348 5740 40404
rect 5796 40348 5806 40404
rect 6738 40348 6748 40404
rect 6804 40348 8092 40404
rect 8148 40348 10556 40404
rect 10612 40348 10622 40404
rect 11414 40348 11452 40404
rect 11508 40348 11518 40404
rect 14354 40348 14364 40404
rect 14420 40348 15596 40404
rect 15652 40348 15662 40404
rect 17714 40348 17724 40404
rect 17780 40348 22540 40404
rect 22596 40348 22606 40404
rect 23426 40348 23436 40404
rect 23492 40348 26572 40404
rect 26628 40348 26638 40404
rect 28354 40348 28364 40404
rect 28420 40348 30156 40404
rect 30212 40348 32172 40404
rect 32228 40348 32238 40404
rect 35298 40348 35308 40404
rect 35364 40348 36316 40404
rect 36372 40348 36382 40404
rect 1698 40236 1708 40292
rect 1764 40236 2492 40292
rect 2548 40236 2558 40292
rect 2818 40236 2828 40292
rect 2884 40236 3388 40292
rect 3444 40236 3482 40292
rect 3602 40236 3612 40292
rect 3668 40236 5628 40292
rect 5684 40236 5694 40292
rect 8194 40236 8204 40292
rect 8260 40236 11788 40292
rect 11844 40236 11854 40292
rect 12898 40236 12908 40292
rect 12964 40236 17556 40292
rect 18498 40236 18508 40292
rect 18564 40236 27916 40292
rect 27972 40236 27982 40292
rect 29474 40236 29484 40292
rect 29540 40236 30828 40292
rect 30884 40236 30894 40292
rect 35186 40236 35196 40292
rect 35252 40236 35868 40292
rect 35924 40236 35934 40292
rect 3388 40180 3444 40236
rect 3388 40124 8092 40180
rect 8148 40124 8158 40180
rect 17500 40068 17556 40236
rect 17714 40124 17724 40180
rect 17780 40124 20636 40180
rect 20692 40124 20702 40180
rect 21522 40124 21532 40180
rect 21588 40124 22652 40180
rect 22708 40124 22718 40180
rect 25666 40124 25676 40180
rect 25732 40124 26348 40180
rect 26404 40124 26414 40180
rect 28242 40124 28252 40180
rect 28308 40124 29372 40180
rect 29428 40124 29438 40180
rect 35522 40124 35532 40180
rect 35588 40124 36428 40180
rect 36484 40124 36494 40180
rect 14690 40012 14700 40068
rect 14756 40012 15036 40068
rect 15092 40012 15102 40068
rect 15362 40012 15372 40068
rect 15428 40012 16604 40068
rect 16660 40012 16670 40068
rect 17500 40012 26124 40068
rect 26180 40012 26190 40068
rect 4466 39956 4476 40012
rect 4532 39956 4580 40012
rect 4636 39956 4684 40012
rect 4740 39956 4750 40012
rect 7746 39788 7756 39844
rect 7812 39788 8204 39844
rect 8260 39788 10332 39844
rect 10388 39788 10398 39844
rect 0 39732 800 39760
rect 15372 39732 15428 40012
rect 16604 39956 16660 40012
rect 35186 39956 35196 40012
rect 35252 39956 35300 40012
rect 35356 39956 35404 40012
rect 35460 39956 35470 40012
rect 16604 39900 19516 39956
rect 19572 39900 19582 39956
rect 28018 39900 28028 39956
rect 28084 39900 28700 39956
rect 28756 39900 29148 39956
rect 29204 39900 29214 39956
rect 15698 39788 15708 39844
rect 15764 39788 16380 39844
rect 16436 39788 20076 39844
rect 20132 39788 20142 39844
rect 21298 39788 21308 39844
rect 21364 39788 22204 39844
rect 22260 39788 22270 39844
rect 26852 39788 30268 39844
rect 30324 39788 30334 39844
rect 26852 39732 26908 39788
rect 0 39676 1708 39732
rect 1764 39676 1774 39732
rect 8306 39676 8316 39732
rect 8372 39676 15428 39732
rect 17378 39676 17388 39732
rect 17444 39676 26908 39732
rect 0 39648 800 39676
rect 1138 39564 1148 39620
rect 1204 39564 2044 39620
rect 2100 39564 2110 39620
rect 2594 39564 2604 39620
rect 2660 39564 3388 39620
rect 3938 39564 3948 39620
rect 4004 39564 5292 39620
rect 5348 39564 6412 39620
rect 6468 39564 6478 39620
rect 7298 39564 7308 39620
rect 7364 39564 7980 39620
rect 8036 39564 8046 39620
rect 10322 39564 10332 39620
rect 10388 39564 10780 39620
rect 10836 39564 12236 39620
rect 12292 39564 12302 39620
rect 26086 39564 26124 39620
rect 26180 39564 26190 39620
rect 26674 39564 26684 39620
rect 26740 39564 28252 39620
rect 28308 39564 28318 39620
rect 29250 39564 29260 39620
rect 29316 39564 30044 39620
rect 30100 39564 30110 39620
rect 3042 39452 3052 39508
rect 3108 39452 3118 39508
rect 3052 39284 3108 39452
rect 3332 39396 3388 39564
rect 5730 39452 5740 39508
rect 5796 39452 12796 39508
rect 12852 39452 12862 39508
rect 14466 39452 14476 39508
rect 14532 39452 14700 39508
rect 14756 39452 18172 39508
rect 18228 39452 18238 39508
rect 23650 39452 23660 39508
rect 23716 39452 23884 39508
rect 23940 39452 23950 39508
rect 26852 39452 27132 39508
rect 27188 39452 27198 39508
rect 32834 39452 32844 39508
rect 32900 39452 33740 39508
rect 33796 39452 33806 39508
rect 26852 39396 26908 39452
rect 3332 39340 3500 39396
rect 3556 39340 3566 39396
rect 10994 39340 11004 39396
rect 11060 39340 11788 39396
rect 11844 39340 11854 39396
rect 14802 39340 14812 39396
rect 14868 39340 19404 39396
rect 19460 39340 20188 39396
rect 20244 39340 24668 39396
rect 24724 39340 24734 39396
rect 25778 39340 25788 39396
rect 25844 39340 26908 39396
rect 27010 39340 27020 39396
rect 27076 39340 31052 39396
rect 31108 39340 31118 39396
rect 3052 39228 3388 39284
rect 3444 39228 3454 39284
rect 10546 39228 10556 39284
rect 10612 39228 13132 39284
rect 13188 39228 13198 39284
rect 14242 39228 14252 39284
rect 14308 39228 18956 39284
rect 19012 39228 19022 39284
rect 20188 39228 24612 39284
rect 24994 39228 25004 39284
rect 25060 39228 25340 39284
rect 25396 39228 25406 39284
rect 25554 39228 25564 39284
rect 25620 39228 26348 39284
rect 26404 39228 26684 39284
rect 26740 39228 26750 39284
rect 31378 39228 31388 39284
rect 31444 39228 33628 39284
rect 33684 39228 33694 39284
rect 19826 39172 19836 39228
rect 19892 39172 19940 39228
rect 19996 39172 20044 39228
rect 20100 39172 20110 39228
rect 11218 39116 11228 39172
rect 11284 39116 15036 39172
rect 15092 39116 15102 39172
rect 20188 39060 20244 39228
rect 24556 39172 24612 39228
rect 50546 39172 50556 39228
rect 50612 39172 50660 39228
rect 50716 39172 50764 39228
rect 50820 39172 50830 39228
rect 24556 39116 28588 39172
rect 28644 39116 28654 39172
rect 3602 39004 3612 39060
rect 3668 39004 5852 39060
rect 5908 39004 5918 39060
rect 7410 39004 7420 39060
rect 7476 39004 7756 39060
rect 7812 39004 7822 39060
rect 13010 39004 13020 39060
rect 13076 39004 14028 39060
rect 14084 39004 14094 39060
rect 14252 39004 20244 39060
rect 20412 39004 24500 39060
rect 25106 39004 25116 39060
rect 25172 39004 25900 39060
rect 25956 39004 25966 39060
rect 14252 38948 14308 39004
rect 3490 38892 3500 38948
rect 3556 38892 5740 38948
rect 5796 38892 5806 38948
rect 6066 38892 6076 38948
rect 6132 38892 14308 38948
rect 15092 38892 16268 38948
rect 16324 38892 16334 38948
rect 18134 38892 18172 38948
rect 18228 38892 18238 38948
rect 6076 38836 6132 38892
rect 15092 38836 15148 38892
rect 20412 38836 20468 39004
rect 24444 38948 24500 39004
rect 22082 38892 22092 38948
rect 22148 38892 24220 38948
rect 24276 38892 24286 38948
rect 24444 38892 27132 38948
rect 27188 38892 27916 38948
rect 27972 38892 27982 38948
rect 35746 38892 35756 38948
rect 35812 38892 38220 38948
rect 38276 38892 38286 38948
rect 3826 38780 3836 38836
rect 3892 38780 4284 38836
rect 4340 38780 6132 38836
rect 6738 38780 6748 38836
rect 6804 38780 10780 38836
rect 10836 38780 10846 38836
rect 12338 38780 12348 38836
rect 12404 38780 15148 38836
rect 15474 38780 15484 38836
rect 15540 38780 16940 38836
rect 16996 38780 17006 38836
rect 18844 38780 20468 38836
rect 20850 38780 20860 38836
rect 20916 38780 21532 38836
rect 21588 38780 21598 38836
rect 21970 38780 21980 38836
rect 22036 38780 26908 38836
rect 26964 38780 26974 38836
rect 18844 38724 18900 38780
rect 6402 38668 6412 38724
rect 6468 38668 8092 38724
rect 8148 38668 8652 38724
rect 8708 38668 8718 38724
rect 15026 38668 15036 38724
rect 15092 38668 18900 38724
rect 22642 38668 22652 38724
rect 22708 38668 23212 38724
rect 23268 38668 23278 38724
rect 23660 38668 25564 38724
rect 25620 38668 25630 38724
rect 25778 38668 25788 38724
rect 25844 38668 25854 38724
rect 26226 38668 26236 38724
rect 26292 38668 27692 38724
rect 27748 38668 27758 38724
rect 34290 38668 34300 38724
rect 34356 38668 34636 38724
rect 34692 38668 34702 38724
rect 35074 38668 35084 38724
rect 35140 38668 36988 38724
rect 37044 38668 37436 38724
rect 37492 38668 37502 38724
rect 9426 38556 9436 38612
rect 9492 38556 23324 38612
rect 23380 38556 23390 38612
rect 23660 38500 23716 38668
rect 25788 38500 25844 38668
rect 13346 38444 13356 38500
rect 13412 38444 23716 38500
rect 24994 38444 25004 38500
rect 25060 38444 25844 38500
rect 31154 38444 31164 38500
rect 31220 38444 32396 38500
rect 32452 38444 32462 38500
rect 4466 38388 4476 38444
rect 4532 38388 4580 38444
rect 4636 38388 4684 38444
rect 4740 38388 4750 38444
rect 35186 38388 35196 38444
rect 35252 38388 35300 38444
rect 35356 38388 35404 38444
rect 35460 38388 35470 38444
rect 2930 38332 2940 38388
rect 2996 38332 3836 38388
rect 3892 38332 3902 38388
rect 11564 38332 14140 38388
rect 14196 38332 14812 38388
rect 14868 38332 14878 38388
rect 15698 38332 15708 38388
rect 15764 38332 16492 38388
rect 16548 38332 16558 38388
rect 19516 38332 22876 38388
rect 22932 38332 22942 38388
rect 24108 38332 27244 38388
rect 27300 38332 27310 38388
rect 4946 38220 4956 38276
rect 5012 38220 9212 38276
rect 9268 38220 9278 38276
rect 9762 38220 9772 38276
rect 9828 38220 11228 38276
rect 11284 38220 11294 38276
rect 11564 38164 11620 38332
rect 19516 38276 19572 38332
rect 24108 38276 24164 38332
rect 12114 38220 12124 38276
rect 12180 38220 13916 38276
rect 13972 38220 14476 38276
rect 14532 38220 14542 38276
rect 16342 38220 16380 38276
rect 16436 38220 16446 38276
rect 16594 38220 16604 38276
rect 16660 38220 19572 38276
rect 19730 38220 19740 38276
rect 19796 38220 21644 38276
rect 21700 38220 21710 38276
rect 21970 38220 21980 38276
rect 22036 38220 24108 38276
rect 24164 38220 24174 38276
rect 26562 38220 26572 38276
rect 26628 38220 26908 38276
rect 28578 38220 28588 38276
rect 28644 38220 37212 38276
rect 37268 38220 37278 38276
rect 37762 38220 37772 38276
rect 37828 38220 39340 38276
rect 39396 38220 39900 38276
rect 39956 38220 39966 38276
rect 26852 38164 26908 38220
rect 3938 38108 3948 38164
rect 4004 38108 11620 38164
rect 12226 38108 12236 38164
rect 12292 38108 12796 38164
rect 12852 38108 20020 38164
rect 22866 38108 22876 38164
rect 22932 38108 25564 38164
rect 25620 38108 25630 38164
rect 26198 38108 26236 38164
rect 26292 38108 26302 38164
rect 26852 38108 28364 38164
rect 28420 38108 28430 38164
rect 30034 38108 30044 38164
rect 30100 38108 31276 38164
rect 31332 38108 34188 38164
rect 34244 38108 34254 38164
rect 19964 38052 20020 38108
rect 4722 37996 4732 38052
rect 4788 37996 8204 38052
rect 8260 37996 8270 38052
rect 10546 37996 10556 38052
rect 10612 37996 15036 38052
rect 15092 37996 15102 38052
rect 15698 37996 15708 38052
rect 15764 37996 16268 38052
rect 16324 37996 16334 38052
rect 17826 37996 17836 38052
rect 17892 37996 18508 38052
rect 18564 37996 18574 38052
rect 19954 37996 19964 38052
rect 20020 37996 20030 38052
rect 23314 37996 23324 38052
rect 23380 37996 26012 38052
rect 26068 37996 26078 38052
rect 30482 37996 30492 38052
rect 30548 37996 31052 38052
rect 31108 37996 32844 38052
rect 32900 37996 32910 38052
rect 36418 37996 36428 38052
rect 36484 37996 38444 38052
rect 38500 37996 38510 38052
rect 0 37940 800 37968
rect 0 37884 1708 37940
rect 1764 37884 1774 37940
rect 13010 37884 13020 37940
rect 13076 37884 15036 37940
rect 15092 37884 16436 37940
rect 17714 37884 17724 37940
rect 17780 37884 19068 37940
rect 19124 37884 19740 37940
rect 19796 37884 19806 37940
rect 24322 37884 24332 37940
rect 24388 37884 24892 37940
rect 24948 37884 24958 37940
rect 28690 37884 28700 37940
rect 28756 37884 30604 37940
rect 30660 37884 30670 37940
rect 32050 37884 32060 37940
rect 32116 37884 33292 37940
rect 33348 37884 33358 37940
rect 0 37856 800 37884
rect 16380 37828 16436 37884
rect 5618 37772 5628 37828
rect 5684 37772 7084 37828
rect 7140 37772 12124 37828
rect 12180 37772 12190 37828
rect 12338 37772 12348 37828
rect 12404 37772 13692 37828
rect 13748 37772 13758 37828
rect 13906 37772 13916 37828
rect 13972 37772 15148 37828
rect 15474 37772 15484 37828
rect 15540 37772 15708 37828
rect 15764 37772 15774 37828
rect 16370 37772 16380 37828
rect 16436 37772 17556 37828
rect 18946 37772 18956 37828
rect 19012 37772 19628 37828
rect 19684 37772 24108 37828
rect 24164 37772 24174 37828
rect 27682 37772 27692 37828
rect 27748 37772 29708 37828
rect 29764 37772 29774 37828
rect 31714 37772 31724 37828
rect 31780 37772 32172 37828
rect 32228 37772 32732 37828
rect 32788 37772 33740 37828
rect 33796 37772 33806 37828
rect 10658 37660 10668 37716
rect 10724 37660 11116 37716
rect 11172 37660 11182 37716
rect 12898 37660 12908 37716
rect 12964 37660 13244 37716
rect 13300 37660 13310 37716
rect 15092 37604 15148 37772
rect 17500 37604 17556 37772
rect 19142 37660 19180 37716
rect 19236 37660 19246 37716
rect 22764 37660 29372 37716
rect 29428 37660 29438 37716
rect 19826 37604 19836 37660
rect 19892 37604 19940 37660
rect 19996 37604 20044 37660
rect 20100 37604 20110 37660
rect 22764 37604 22820 37660
rect 50546 37604 50556 37660
rect 50612 37604 50660 37660
rect 50716 37604 50764 37660
rect 50820 37604 50830 37660
rect 3602 37548 3612 37604
rect 3668 37548 3948 37604
rect 4004 37548 4014 37604
rect 13906 37548 13916 37604
rect 13972 37548 14364 37604
rect 14420 37548 14430 37604
rect 15092 37548 16492 37604
rect 16548 37548 16558 37604
rect 17490 37548 17500 37604
rect 17556 37548 17566 37604
rect 18246 37548 18284 37604
rect 18340 37548 18350 37604
rect 21074 37548 21084 37604
rect 21140 37548 21980 37604
rect 22036 37548 22046 37604
rect 22754 37548 22764 37604
rect 22820 37548 22830 37604
rect 24546 37548 24556 37604
rect 24612 37548 25676 37604
rect 25732 37548 25742 37604
rect 1922 37436 1932 37492
rect 1988 37436 2604 37492
rect 2660 37436 2670 37492
rect 2818 37436 2828 37492
rect 2884 37436 17276 37492
rect 17332 37436 17342 37492
rect 18386 37436 18396 37492
rect 18452 37436 19180 37492
rect 19236 37436 19246 37492
rect 19394 37436 19404 37492
rect 19460 37436 21420 37492
rect 21476 37436 21486 37492
rect 21644 37436 25228 37492
rect 25284 37436 25294 37492
rect 26758 37436 26796 37492
rect 26852 37436 26862 37492
rect 29586 37436 29596 37492
rect 29652 37436 31500 37492
rect 31556 37436 31724 37492
rect 31780 37436 32060 37492
rect 32116 37436 32126 37492
rect 21644 37380 21700 37436
rect 8978 37324 8988 37380
rect 9044 37324 9212 37380
rect 9268 37324 9278 37380
rect 11890 37324 11900 37380
rect 11956 37324 12572 37380
rect 12628 37324 12638 37380
rect 15138 37324 15148 37380
rect 15204 37324 16156 37380
rect 16212 37324 16222 37380
rect 16482 37324 16492 37380
rect 16548 37324 18284 37380
rect 18340 37324 21700 37380
rect 21970 37324 21980 37380
rect 22036 37324 22764 37380
rect 22820 37324 22830 37380
rect 24658 37324 24668 37380
rect 24724 37324 26236 37380
rect 26292 37324 29036 37380
rect 29092 37324 29484 37380
rect 29540 37324 29550 37380
rect 38098 37324 38108 37380
rect 38164 37324 39564 37380
rect 39620 37324 39630 37380
rect 3602 37212 3612 37268
rect 3668 37212 10108 37268
rect 10164 37212 10174 37268
rect 12870 37212 12908 37268
rect 12964 37212 12974 37268
rect 13682 37212 13692 37268
rect 13748 37212 16100 37268
rect 16258 37212 16268 37268
rect 16324 37212 17388 37268
rect 17444 37212 17454 37268
rect 17826 37212 17836 37268
rect 17892 37212 18396 37268
rect 18452 37212 18462 37268
rect 21186 37212 21196 37268
rect 21252 37212 22540 37268
rect 22596 37212 22606 37268
rect 25442 37212 25452 37268
rect 25508 37212 26572 37268
rect 26628 37212 27468 37268
rect 27524 37212 27534 37268
rect 27692 37212 28028 37268
rect 28084 37212 28094 37268
rect 32386 37212 32396 37268
rect 32452 37212 34188 37268
rect 34244 37212 35644 37268
rect 35700 37212 35710 37268
rect 1698 37100 1708 37156
rect 1764 37100 3164 37156
rect 3220 37100 3230 37156
rect 7410 37100 7420 37156
rect 7476 37100 8428 37156
rect 8484 37100 15988 37156
rect 8978 36988 8988 37044
rect 9044 36988 9660 37044
rect 9716 36988 9726 37044
rect 11106 36988 11116 37044
rect 11172 36988 12124 37044
rect 12180 36988 13356 37044
rect 13412 36988 13422 37044
rect 13570 36988 13580 37044
rect 13636 36988 14028 37044
rect 14084 36988 14094 37044
rect 15932 36932 15988 37100
rect 16044 37044 16100 37212
rect 27692 37156 27748 37212
rect 18610 37100 18620 37156
rect 18676 37100 21084 37156
rect 21140 37100 21150 37156
rect 21410 37100 21420 37156
rect 21476 37100 25228 37156
rect 25284 37100 25294 37156
rect 25554 37100 25564 37156
rect 25620 37100 27748 37156
rect 27906 37100 27916 37156
rect 27972 37100 28588 37156
rect 28644 37100 29036 37156
rect 29092 37100 29102 37156
rect 30034 37100 30044 37156
rect 30100 37100 31948 37156
rect 32004 37100 32014 37156
rect 37986 37100 37996 37156
rect 38052 37100 38668 37156
rect 38724 37100 38734 37156
rect 16044 36988 21532 37044
rect 21588 36988 22988 37044
rect 23044 36988 23054 37044
rect 25778 36988 25788 37044
rect 25844 36988 30492 37044
rect 30548 36988 30558 37044
rect 15932 36876 19180 36932
rect 19236 36876 19404 36932
rect 19460 36876 20412 36932
rect 20468 36876 20748 36932
rect 20804 36876 23212 36932
rect 23268 36876 23278 36932
rect 23426 36876 23436 36932
rect 23492 36876 26124 36932
rect 26180 36876 26190 36932
rect 26898 36876 26908 36932
rect 26964 36876 27356 36932
rect 27412 36876 27916 36932
rect 27972 36876 27982 36932
rect 4466 36820 4476 36876
rect 4532 36820 4580 36876
rect 4636 36820 4684 36876
rect 4740 36820 4750 36876
rect 15026 36764 15036 36820
rect 15092 36764 18396 36820
rect 18452 36764 18462 36820
rect 14130 36652 14140 36708
rect 14196 36652 14924 36708
rect 14980 36652 14990 36708
rect 18050 36652 18060 36708
rect 18116 36652 18508 36708
rect 18564 36652 18574 36708
rect 3126 36540 3164 36596
rect 3220 36540 3230 36596
rect 11442 36540 11452 36596
rect 11508 36540 19180 36596
rect 19236 36540 19246 36596
rect 19842 36540 19852 36596
rect 19908 36540 21868 36596
rect 21924 36540 21934 36596
rect 23212 36484 23268 36876
rect 35186 36820 35196 36876
rect 35252 36820 35300 36876
rect 35356 36820 35404 36876
rect 35460 36820 35470 36876
rect 26562 36764 26572 36820
rect 26628 36764 29932 36820
rect 29988 36764 29998 36820
rect 25330 36652 25340 36708
rect 25396 36652 26012 36708
rect 26068 36652 26908 36708
rect 26852 36596 26908 36652
rect 26852 36540 27580 36596
rect 27636 36540 27646 36596
rect 2034 36428 2044 36484
rect 2100 36428 2716 36484
rect 2772 36428 2782 36484
rect 2940 36428 3276 36484
rect 3332 36428 3342 36484
rect 12898 36428 12908 36484
rect 12964 36428 13804 36484
rect 13860 36428 13870 36484
rect 14354 36428 14364 36484
rect 14420 36428 17948 36484
rect 18004 36428 20860 36484
rect 20916 36428 20926 36484
rect 23212 36428 25340 36484
rect 25396 36428 25406 36484
rect 26852 36428 28476 36484
rect 28532 36428 28542 36484
rect 33170 36428 33180 36484
rect 33236 36428 37996 36484
rect 38052 36428 38062 36484
rect 2940 36372 2996 36428
rect 26852 36372 26908 36428
rect 1362 36316 1372 36372
rect 1428 36316 1932 36372
rect 1988 36316 1998 36372
rect 2370 36316 2380 36372
rect 2436 36316 2996 36372
rect 5618 36316 5628 36372
rect 5684 36316 5964 36372
rect 6020 36316 6748 36372
rect 6804 36316 6814 36372
rect 17490 36316 17500 36372
rect 17556 36316 21924 36372
rect 24210 36316 24220 36372
rect 24276 36316 26908 36372
rect 28018 36316 28028 36372
rect 28084 36316 28364 36372
rect 28420 36316 28430 36372
rect 0 36148 800 36176
rect 0 36092 1708 36148
rect 1764 36092 1774 36148
rect 0 36064 800 36092
rect 1932 35924 1988 36316
rect 21868 36260 21924 36316
rect 10322 36204 10332 36260
rect 10388 36204 10556 36260
rect 10612 36204 11116 36260
rect 11172 36204 12572 36260
rect 12628 36204 12638 36260
rect 14914 36204 14924 36260
rect 14980 36204 16380 36260
rect 16436 36204 17836 36260
rect 17892 36204 17902 36260
rect 18358 36204 18396 36260
rect 18452 36204 18462 36260
rect 18610 36204 18620 36260
rect 18676 36204 18956 36260
rect 19012 36204 19022 36260
rect 20290 36204 20300 36260
rect 20356 36204 20366 36260
rect 21858 36204 21868 36260
rect 21924 36204 21934 36260
rect 22092 36204 28476 36260
rect 28532 36204 29260 36260
rect 29316 36204 29326 36260
rect 29698 36204 29708 36260
rect 29764 36204 29774 36260
rect 33842 36204 33852 36260
rect 33908 36204 33918 36260
rect 38994 36204 39004 36260
rect 39060 36204 40124 36260
rect 40180 36204 40190 36260
rect 20300 36148 20356 36204
rect 22092 36148 22148 36204
rect 2790 36092 2828 36148
rect 2884 36092 2894 36148
rect 7746 36092 7756 36148
rect 7812 36092 12012 36148
rect 12068 36092 12078 36148
rect 13122 36092 13132 36148
rect 13188 36092 13692 36148
rect 13748 36092 13758 36148
rect 15138 36092 15148 36148
rect 15204 36092 17724 36148
rect 17780 36092 17790 36148
rect 18162 36092 18172 36148
rect 18228 36092 18284 36148
rect 18340 36092 18350 36148
rect 19170 36092 19180 36148
rect 19236 36092 19292 36148
rect 19348 36092 19358 36148
rect 20300 36092 22148 36148
rect 22530 36092 22540 36148
rect 22596 36092 26908 36148
rect 27990 36092 28028 36148
rect 28084 36092 28094 36148
rect 19826 36036 19836 36092
rect 19892 36036 19940 36092
rect 19996 36036 20044 36092
rect 20100 36036 20110 36092
rect 26852 36036 26908 36092
rect 29708 36036 29764 36204
rect 4274 35980 4284 36036
rect 4340 35980 17780 36036
rect 1932 35868 4620 35924
rect 4676 35868 4686 35924
rect 6300 35868 10108 35924
rect 10164 35868 10174 35924
rect 12002 35868 12012 35924
rect 12068 35868 13916 35924
rect 13972 35868 13982 35924
rect 15026 35868 15036 35924
rect 15092 35868 16044 35924
rect 16100 35868 16110 35924
rect 1026 35756 1036 35812
rect 1092 35756 2716 35812
rect 2772 35756 2782 35812
rect 6300 35700 6356 35868
rect 17724 35812 17780 35980
rect 20636 35980 20972 36036
rect 21028 35980 21038 36036
rect 26852 35980 30940 36036
rect 30996 35980 31006 36036
rect 20636 35924 20692 35980
rect 33852 35924 33908 36204
rect 50546 36036 50556 36092
rect 50612 36036 50660 36092
rect 50716 36036 50764 36092
rect 50820 36036 50830 36092
rect 38434 35980 38444 36036
rect 38500 35980 40348 36036
rect 40404 35980 40908 36036
rect 40964 35980 40974 36036
rect 19842 35868 19852 35924
rect 19908 35868 20692 35924
rect 20850 35868 20860 35924
rect 20916 35868 22876 35924
rect 22932 35868 22942 35924
rect 23538 35868 23548 35924
rect 23604 35868 25676 35924
rect 25732 35868 33908 35924
rect 34402 35868 34412 35924
rect 34468 35868 35532 35924
rect 35588 35868 36428 35924
rect 36484 35868 39228 35924
rect 39284 35868 39294 35924
rect 8978 35756 8988 35812
rect 9044 35756 15148 35812
rect 17714 35756 17724 35812
rect 17780 35756 17790 35812
rect 18806 35756 18844 35812
rect 18900 35756 18910 35812
rect 19282 35756 19292 35812
rect 19348 35756 24332 35812
rect 24388 35756 25340 35812
rect 25396 35756 25406 35812
rect 35634 35756 35644 35812
rect 35700 35756 37436 35812
rect 37492 35756 37502 35812
rect 15092 35700 15148 35756
rect 2594 35644 2604 35700
rect 2660 35644 6356 35700
rect 8530 35644 8540 35700
rect 8596 35644 10444 35700
rect 10500 35644 10510 35700
rect 12002 35644 12012 35700
rect 12068 35644 13468 35700
rect 13524 35644 13534 35700
rect 15092 35644 20300 35700
rect 20356 35644 20366 35700
rect 27766 35644 27804 35700
rect 27860 35644 28812 35700
rect 28868 35644 31724 35700
rect 31780 35644 31790 35700
rect 32274 35644 32284 35700
rect 32340 35644 34972 35700
rect 35028 35644 35038 35700
rect 36194 35644 36204 35700
rect 36260 35644 37100 35700
rect 37156 35644 39004 35700
rect 39060 35644 39070 35700
rect 12012 35588 12068 35644
rect 2818 35532 2828 35588
rect 2884 35532 3052 35588
rect 3108 35532 3118 35588
rect 3490 35532 3500 35588
rect 3556 35532 4284 35588
rect 4340 35532 4350 35588
rect 5394 35532 5404 35588
rect 5460 35532 12068 35588
rect 15362 35532 15372 35588
rect 15428 35532 16268 35588
rect 16324 35532 16334 35588
rect 20066 35532 20076 35588
rect 20132 35532 21420 35588
rect 21476 35532 21486 35588
rect 21634 35532 21644 35588
rect 21700 35532 27132 35588
rect 27188 35532 27198 35588
rect 39666 35532 39676 35588
rect 39732 35532 41356 35588
rect 41412 35532 41422 35588
rect 3938 35420 3948 35476
rect 4004 35420 9772 35476
rect 9828 35420 9838 35476
rect 10210 35420 10220 35476
rect 10276 35420 10286 35476
rect 10546 35420 10556 35476
rect 10612 35420 10780 35476
rect 10836 35420 10846 35476
rect 13132 35420 14140 35476
rect 14196 35420 18620 35476
rect 18676 35420 20860 35476
rect 20916 35420 26684 35476
rect 26740 35420 27580 35476
rect 27636 35420 28476 35476
rect 28532 35420 28542 35476
rect 34738 35420 34748 35476
rect 34804 35420 36316 35476
rect 36372 35420 36382 35476
rect 4834 35308 4844 35364
rect 4900 35308 5740 35364
rect 5796 35308 5806 35364
rect 8194 35308 8204 35364
rect 8260 35308 9884 35364
rect 9940 35308 9950 35364
rect 10220 35308 10276 35420
rect 13132 35364 13188 35420
rect 10434 35308 10444 35364
rect 10500 35308 13188 35364
rect 14914 35308 14924 35364
rect 14980 35308 15372 35364
rect 15428 35308 15438 35364
rect 17042 35308 17052 35364
rect 17108 35308 18956 35364
rect 19012 35308 19022 35364
rect 19954 35308 19964 35364
rect 20020 35308 20300 35364
rect 20356 35308 20366 35364
rect 20962 35308 20972 35364
rect 21028 35308 22876 35364
rect 22932 35308 22942 35364
rect 23874 35308 23884 35364
rect 23940 35308 26012 35364
rect 26068 35308 26078 35364
rect 27122 35308 27132 35364
rect 27188 35308 27804 35364
rect 27860 35308 27870 35364
rect 36418 35308 36428 35364
rect 36484 35308 39116 35364
rect 39172 35308 39182 35364
rect 4466 35252 4476 35308
rect 4532 35252 4580 35308
rect 4636 35252 4684 35308
rect 4740 35252 4750 35308
rect 10210 35252 10220 35308
rect 10276 35252 10286 35308
rect 35186 35252 35196 35308
rect 35252 35252 35300 35308
rect 35356 35252 35404 35308
rect 35460 35252 35470 35308
rect 18806 35196 18844 35252
rect 18900 35196 18910 35252
rect 19170 35196 19180 35252
rect 19236 35196 23772 35252
rect 23828 35196 25340 35252
rect 25396 35196 25406 35252
rect 26226 35196 26236 35252
rect 26292 35196 29372 35252
rect 29428 35196 29438 35252
rect 29810 35196 29820 35252
rect 29876 35196 30940 35252
rect 30996 35196 33404 35252
rect 33460 35196 33470 35252
rect 6290 35084 6300 35140
rect 6356 35084 11564 35140
rect 11620 35084 12236 35140
rect 12292 35084 12302 35140
rect 18470 35084 18508 35140
rect 18564 35084 18574 35140
rect 19366 35084 19404 35140
rect 19460 35084 19470 35140
rect 27010 35084 27020 35140
rect 27076 35084 29260 35140
rect 29316 35084 29326 35140
rect 31602 35084 31612 35140
rect 31668 35084 33180 35140
rect 33236 35084 35532 35140
rect 35588 35084 35598 35140
rect 38658 35084 38668 35140
rect 38724 35084 39340 35140
rect 39396 35084 39406 35140
rect 9874 34972 9884 35028
rect 9940 34972 10444 35028
rect 10500 34972 14700 35028
rect 14756 34972 14766 35028
rect 15922 34972 15932 35028
rect 15988 34972 24108 35028
rect 24164 34972 24668 35028
rect 24724 34972 25732 35028
rect 26450 34972 26460 35028
rect 26516 34972 27132 35028
rect 27188 34972 27198 35028
rect 28578 34972 28588 35028
rect 28644 34972 29708 35028
rect 29764 34972 29774 35028
rect 25676 34916 25732 34972
rect 2146 34860 2156 34916
rect 2212 34860 2604 34916
rect 2660 34860 2670 34916
rect 12562 34860 12572 34916
rect 12628 34860 13468 34916
rect 13524 34860 13534 34916
rect 14438 34860 14476 34916
rect 14532 34860 14542 34916
rect 16902 34860 16940 34916
rect 16996 34860 17006 34916
rect 18498 34860 18508 34916
rect 18564 34860 25452 34916
rect 25508 34860 25518 34916
rect 25676 34860 26684 34916
rect 26740 34860 26750 34916
rect 36866 34860 36876 34916
rect 36932 34860 38556 34916
rect 38612 34860 38622 34916
rect 11554 34748 11564 34804
rect 11620 34748 16828 34804
rect 16884 34748 16894 34804
rect 18274 34748 18284 34804
rect 18340 34748 18844 34804
rect 18900 34748 22764 34804
rect 22820 34748 22830 34804
rect 31714 34748 31724 34804
rect 31780 34748 35588 34804
rect 36306 34748 36316 34804
rect 36372 34748 37100 34804
rect 37156 34748 37660 34804
rect 37716 34748 41468 34804
rect 41524 34748 41534 34804
rect 35532 34692 35588 34748
rect 2930 34636 2940 34692
rect 2996 34636 3164 34692
rect 3220 34636 5292 34692
rect 5348 34636 5358 34692
rect 6178 34636 6188 34692
rect 6244 34636 7868 34692
rect 7924 34636 7934 34692
rect 11330 34636 11340 34692
rect 11396 34636 13580 34692
rect 13636 34636 13646 34692
rect 14354 34636 14364 34692
rect 14420 34636 14700 34692
rect 14756 34636 14766 34692
rect 19058 34636 19068 34692
rect 19124 34636 19740 34692
rect 19796 34636 22652 34692
rect 22708 34636 22718 34692
rect 28018 34636 28028 34692
rect 28084 34636 28700 34692
rect 28756 34636 30380 34692
rect 30436 34636 30446 34692
rect 30706 34636 30716 34692
rect 30772 34636 35308 34692
rect 35364 34636 35374 34692
rect 35532 34636 37212 34692
rect 37268 34636 37278 34692
rect 2818 34524 2828 34580
rect 2884 34524 3164 34580
rect 3220 34524 3230 34580
rect 9650 34524 9660 34580
rect 9716 34524 13916 34580
rect 13972 34524 15148 34580
rect 21858 34524 21868 34580
rect 21924 34524 23772 34580
rect 23828 34524 23838 34580
rect 15092 34468 15148 34524
rect 19826 34468 19836 34524
rect 19892 34468 19940 34524
rect 19996 34468 20044 34524
rect 20100 34468 20110 34524
rect 28028 34468 28084 34636
rect 50546 34468 50556 34524
rect 50612 34468 50660 34524
rect 50716 34468 50764 34524
rect 50820 34468 50830 34524
rect 8082 34412 8092 34468
rect 8148 34412 12012 34468
rect 12068 34412 12078 34468
rect 14242 34412 14252 34468
rect 14308 34412 14364 34468
rect 14420 34412 14430 34468
rect 14802 34412 14812 34468
rect 14868 34412 14878 34468
rect 15092 34412 17948 34468
rect 18004 34412 19292 34468
rect 19348 34412 19358 34468
rect 20962 34412 20972 34468
rect 21028 34412 28084 34468
rect 0 34356 800 34384
rect 14812 34356 14868 34412
rect 0 34300 1708 34356
rect 1764 34300 1774 34356
rect 4386 34300 4396 34356
rect 4452 34300 5404 34356
rect 5460 34300 5470 34356
rect 6626 34300 6636 34356
rect 6692 34300 8540 34356
rect 8596 34300 8606 34356
rect 9650 34300 9660 34356
rect 9716 34300 10108 34356
rect 10164 34300 10174 34356
rect 11666 34300 11676 34356
rect 11732 34300 11742 34356
rect 14812 34300 15036 34356
rect 15092 34300 17332 34356
rect 17574 34300 17612 34356
rect 17668 34300 17678 34356
rect 21634 34300 21644 34356
rect 21700 34300 28252 34356
rect 28308 34300 29260 34356
rect 29316 34300 29326 34356
rect 0 34272 800 34300
rect 11676 34244 11732 34300
rect 2034 34188 2044 34244
rect 2100 34188 6524 34244
rect 6580 34188 6590 34244
rect 10546 34188 10556 34244
rect 10612 34188 11116 34244
rect 11172 34188 11182 34244
rect 11676 34188 17052 34244
rect 17108 34188 17118 34244
rect 17276 34132 17332 34300
rect 17490 34188 17500 34244
rect 17556 34188 26236 34244
rect 26292 34188 26302 34244
rect 15586 34076 15596 34132
rect 15652 34076 16716 34132
rect 16772 34076 16782 34132
rect 17276 34076 19068 34132
rect 19124 34076 19134 34132
rect 19282 34076 19292 34132
rect 19348 34076 19516 34132
rect 19572 34076 20972 34132
rect 21028 34076 21038 34132
rect 21298 34076 21308 34132
rect 21364 34076 21868 34132
rect 21924 34076 23996 34132
rect 24052 34076 24062 34132
rect 26786 34076 26796 34132
rect 26852 34076 27020 34132
rect 27076 34076 27086 34132
rect 35410 34076 35420 34132
rect 35476 34076 36092 34132
rect 36148 34076 36158 34132
rect 36418 34076 36428 34132
rect 36484 34076 39564 34132
rect 39620 34076 40124 34132
rect 40180 34076 40190 34132
rect 7522 33964 7532 34020
rect 7588 33964 8204 34020
rect 8260 33964 8270 34020
rect 10098 33964 10108 34020
rect 10164 33964 10668 34020
rect 10724 33964 10734 34020
rect 12002 33964 12012 34020
rect 12068 33964 12908 34020
rect 12964 33964 12974 34020
rect 14914 33964 14924 34020
rect 14980 33964 17612 34020
rect 17668 33964 17678 34020
rect 18050 33964 18060 34020
rect 18116 33964 19180 34020
rect 19236 33964 19246 34020
rect 20262 33964 20300 34020
rect 20356 33964 20366 34020
rect 21858 33964 21868 34020
rect 21924 33964 30268 34020
rect 30324 33964 30334 34020
rect 14690 33852 14700 33908
rect 14756 33852 17724 33908
rect 17780 33852 18396 33908
rect 18452 33852 18462 33908
rect 22642 33852 22652 33908
rect 22708 33852 23772 33908
rect 23828 33852 23838 33908
rect 26450 33852 26460 33908
rect 26516 33852 27580 33908
rect 27636 33852 27646 33908
rect 11106 33740 11116 33796
rect 11172 33740 16436 33796
rect 16930 33740 16940 33796
rect 16996 33740 17948 33796
rect 18004 33740 21196 33796
rect 21252 33740 21262 33796
rect 4466 33684 4476 33740
rect 4532 33684 4580 33740
rect 4636 33684 4684 33740
rect 4740 33684 4750 33740
rect 13234 33628 13244 33684
rect 13300 33628 14028 33684
rect 14084 33628 14094 33684
rect 3042 33516 3052 33572
rect 3108 33516 4620 33572
rect 4676 33516 4686 33572
rect 6598 33516 6636 33572
rect 6692 33516 6702 33572
rect 14242 33516 14252 33572
rect 14308 33516 14588 33572
rect 14644 33516 14654 33572
rect 16380 33460 16436 33740
rect 35186 33684 35196 33740
rect 35252 33684 35300 33740
rect 35356 33684 35404 33740
rect 35460 33684 35470 33740
rect 16594 33628 16604 33684
rect 16660 33628 16670 33684
rect 17042 33628 17052 33684
rect 17108 33628 20860 33684
rect 20916 33628 21644 33684
rect 21700 33628 21710 33684
rect 25330 33628 25340 33684
rect 25396 33628 27244 33684
rect 27300 33628 27804 33684
rect 27860 33628 27870 33684
rect 36082 33628 36092 33684
rect 36148 33628 37324 33684
rect 37380 33628 38220 33684
rect 38276 33628 38286 33684
rect 38882 33628 38892 33684
rect 38948 33628 38958 33684
rect 16604 33572 16660 33628
rect 38892 33572 38948 33628
rect 16604 33516 17388 33572
rect 17444 33516 17454 33572
rect 19058 33516 19068 33572
rect 19124 33516 25508 33572
rect 31378 33516 31388 33572
rect 31444 33516 32172 33572
rect 32228 33516 32238 33572
rect 32386 33516 32396 33572
rect 32452 33516 33292 33572
rect 33348 33516 34300 33572
rect 34356 33516 34366 33572
rect 38892 33516 39676 33572
rect 39732 33516 39742 33572
rect 9202 33404 9212 33460
rect 9268 33404 9660 33460
rect 9716 33404 10444 33460
rect 10500 33404 10780 33460
rect 10836 33404 10846 33460
rect 13010 33404 13020 33460
rect 13076 33404 13244 33460
rect 13300 33404 15484 33460
rect 15540 33404 15550 33460
rect 16380 33404 17556 33460
rect 18274 33404 18284 33460
rect 18340 33404 19180 33460
rect 19236 33404 19246 33460
rect 22082 33404 22092 33460
rect 22148 33404 22988 33460
rect 23044 33404 23054 33460
rect 23314 33404 23324 33460
rect 23380 33404 25228 33460
rect 25284 33404 25294 33460
rect 17500 33348 17556 33404
rect 25452 33348 25508 33516
rect 38892 33460 38948 33516
rect 33170 33404 33180 33460
rect 33236 33404 38948 33460
rect 2258 33292 2268 33348
rect 2324 33292 2828 33348
rect 2884 33292 2894 33348
rect 5058 33292 5068 33348
rect 5124 33292 5964 33348
rect 6020 33292 6030 33348
rect 8642 33292 8652 33348
rect 8708 33292 17332 33348
rect 17490 33292 17500 33348
rect 17556 33292 19292 33348
rect 19348 33292 19358 33348
rect 22306 33292 22316 33348
rect 22372 33292 23436 33348
rect 23492 33292 25116 33348
rect 25172 33292 25182 33348
rect 25452 33292 26908 33348
rect 27010 33292 27020 33348
rect 27076 33292 27356 33348
rect 27412 33292 27422 33348
rect 28018 33292 28028 33348
rect 28084 33292 28812 33348
rect 28868 33292 28878 33348
rect 37090 33292 37100 33348
rect 37156 33292 39452 33348
rect 39508 33292 40908 33348
rect 40964 33292 40974 33348
rect 17276 33236 17332 33292
rect 1698 33180 1708 33236
rect 1764 33180 2492 33236
rect 2548 33180 2558 33236
rect 3154 33180 3164 33236
rect 3220 33180 4284 33236
rect 4340 33180 5180 33236
rect 5236 33180 5246 33236
rect 7074 33180 7084 33236
rect 7140 33180 14028 33236
rect 14084 33180 15932 33236
rect 15988 33180 15998 33236
rect 16146 33180 16156 33236
rect 16212 33180 16380 33236
rect 16436 33180 16446 33236
rect 17276 33180 18284 33236
rect 18340 33180 20636 33236
rect 20692 33180 20702 33236
rect 22082 33180 22092 33236
rect 22148 33180 25340 33236
rect 25396 33180 25406 33236
rect 26852 33124 26908 33292
rect 28242 33180 28252 33236
rect 28308 33180 29260 33236
rect 29316 33180 29326 33236
rect 33842 33180 33852 33236
rect 33908 33180 35644 33236
rect 35700 33180 35710 33236
rect 2034 33068 2044 33124
rect 2100 33068 3612 33124
rect 3668 33068 3678 33124
rect 10658 33068 10668 33124
rect 10724 33068 13020 33124
rect 13076 33068 13086 33124
rect 15026 33068 15036 33124
rect 15092 33068 16940 33124
rect 16996 33068 17006 33124
rect 17154 33068 17164 33124
rect 17220 33068 18620 33124
rect 18676 33068 18956 33124
rect 19012 33068 19022 33124
rect 19394 33068 19404 33124
rect 19460 33068 19516 33124
rect 19572 33068 19964 33124
rect 20020 33068 20030 33124
rect 20850 33068 20860 33124
rect 20916 33068 23212 33124
rect 23268 33068 23278 33124
rect 26852 33068 27692 33124
rect 27748 33068 29148 33124
rect 29204 33068 29214 33124
rect 37202 33068 37212 33124
rect 37268 33068 38668 33124
rect 38724 33068 38734 33124
rect 7634 32956 7644 33012
rect 7700 32956 17948 33012
rect 18004 32956 18014 33012
rect 18162 32956 18172 33012
rect 18228 32956 18284 33012
rect 18340 32956 18350 33012
rect 20290 32956 20300 33012
rect 20356 32956 22764 33012
rect 22820 32956 24220 33012
rect 24276 32956 24286 33012
rect 24434 32956 24444 33012
rect 24500 32956 33852 33012
rect 33908 32956 33918 33012
rect 15036 32900 15092 32956
rect 19826 32900 19836 32956
rect 19892 32900 19940 32956
rect 19996 32900 20044 32956
rect 20100 32900 20110 32956
rect 50546 32900 50556 32956
rect 50612 32900 50660 32956
rect 50716 32900 50764 32956
rect 50820 32900 50830 32956
rect 8866 32844 8876 32900
rect 8932 32844 9660 32900
rect 9716 32844 9726 32900
rect 15026 32844 15036 32900
rect 15092 32844 15102 32900
rect 20178 32844 20188 32900
rect 20244 32844 20282 32900
rect 34738 32844 34748 32900
rect 34804 32844 34972 32900
rect 35028 32844 36428 32900
rect 36484 32844 39116 32900
rect 39172 32844 39182 32900
rect 11890 32732 11900 32788
rect 11956 32732 21644 32788
rect 21700 32732 23436 32788
rect 23492 32732 27580 32788
rect 27636 32732 28028 32788
rect 28084 32732 28094 32788
rect 32162 32732 32172 32788
rect 32228 32732 37660 32788
rect 37716 32732 37726 32788
rect 10882 32620 10892 32676
rect 10948 32620 13916 32676
rect 13972 32620 14252 32676
rect 14308 32620 14318 32676
rect 14578 32620 14588 32676
rect 14644 32620 19516 32676
rect 19572 32620 19582 32676
rect 20850 32620 20860 32676
rect 20916 32620 23100 32676
rect 23156 32620 23166 32676
rect 26562 32620 26572 32676
rect 26628 32620 27020 32676
rect 27076 32620 28364 32676
rect 28420 32620 28430 32676
rect 33394 32620 33404 32676
rect 33460 32620 34524 32676
rect 34580 32620 37324 32676
rect 37380 32620 37390 32676
rect 0 32564 800 32592
rect 14252 32564 14308 32620
rect 0 32508 1708 32564
rect 1764 32508 1774 32564
rect 3332 32508 4956 32564
rect 5012 32508 7308 32564
rect 7364 32508 7374 32564
rect 10406 32508 10444 32564
rect 10500 32508 10510 32564
rect 13122 32508 13132 32564
rect 13188 32508 13580 32564
rect 13636 32508 13646 32564
rect 14252 32508 16828 32564
rect 16884 32508 17724 32564
rect 17780 32508 17790 32564
rect 17938 32508 17948 32564
rect 18004 32508 22540 32564
rect 22596 32508 22606 32564
rect 22978 32508 22988 32564
rect 23044 32508 25340 32564
rect 25396 32508 25406 32564
rect 25564 32508 27692 32564
rect 27748 32508 27758 32564
rect 28914 32508 28924 32564
rect 28980 32508 29484 32564
rect 29540 32508 29550 32564
rect 34178 32508 34188 32564
rect 34244 32508 34748 32564
rect 34804 32508 35196 32564
rect 35252 32508 35262 32564
rect 0 32480 800 32508
rect 3332 32452 3388 32508
rect 22540 32452 22596 32508
rect 25564 32452 25620 32508
rect 1250 32396 1260 32452
rect 1316 32396 3388 32452
rect 16482 32396 16492 32452
rect 16548 32396 18060 32452
rect 18116 32396 19964 32452
rect 20020 32396 21420 32452
rect 21476 32396 21486 32452
rect 22540 32396 24668 32452
rect 24724 32396 25564 32452
rect 25620 32396 25630 32452
rect 6626 32284 6636 32340
rect 6692 32284 11004 32340
rect 11060 32284 11070 32340
rect 12450 32284 12460 32340
rect 12516 32284 12796 32340
rect 12852 32284 16604 32340
rect 16660 32284 16670 32340
rect 16818 32284 16828 32340
rect 16884 32284 21084 32340
rect 21140 32284 21150 32340
rect 10098 32172 10108 32228
rect 10164 32172 22092 32228
rect 22148 32172 23436 32228
rect 23492 32172 23502 32228
rect 4466 32116 4476 32172
rect 4532 32116 4580 32172
rect 4636 32116 4684 32172
rect 4740 32116 4750 32172
rect 35186 32116 35196 32172
rect 35252 32116 35300 32172
rect 35356 32116 35404 32172
rect 35460 32116 35470 32172
rect 3714 32060 3724 32116
rect 3780 32060 4060 32116
rect 4116 32060 4126 32116
rect 12450 32060 12460 32116
rect 12516 32060 13356 32116
rect 13412 32060 13422 32116
rect 19170 32060 19180 32116
rect 19236 32060 19852 32116
rect 19908 32060 19918 32116
rect 5618 31948 5628 32004
rect 5684 31948 7084 32004
rect 7140 31948 7150 32004
rect 13122 31948 13132 32004
rect 13188 31948 14028 32004
rect 14084 31948 15260 32004
rect 15316 31948 15326 32004
rect 16146 31948 16156 32004
rect 16212 31948 16716 32004
rect 16772 31948 16782 32004
rect 17042 31948 17052 32004
rect 17108 31948 17612 32004
rect 17668 31948 17678 32004
rect 18834 31948 18844 32004
rect 18900 31948 24332 32004
rect 24388 31948 24398 32004
rect 2930 31836 2940 31892
rect 2996 31836 3612 31892
rect 3668 31836 3678 31892
rect 9090 31836 9100 31892
rect 9156 31836 9548 31892
rect 9604 31836 13356 31892
rect 13412 31836 13422 31892
rect 20066 31836 20076 31892
rect 20132 31836 20300 31892
rect 20356 31836 20366 31892
rect 20850 31836 20860 31892
rect 20916 31836 22988 31892
rect 23044 31836 23054 31892
rect 3378 31724 3388 31780
rect 3444 31724 3724 31780
rect 3780 31724 3790 31780
rect 13906 31724 13916 31780
rect 13972 31724 14812 31780
rect 14868 31724 14878 31780
rect 15092 31724 16604 31780
rect 16660 31724 16670 31780
rect 18498 31724 18508 31780
rect 18564 31724 20188 31780
rect 20244 31724 21868 31780
rect 21924 31724 22316 31780
rect 22372 31724 22382 31780
rect 22530 31724 22540 31780
rect 22596 31724 22764 31780
rect 22820 31724 23660 31780
rect 23716 31724 24444 31780
rect 24500 31724 24510 31780
rect 15092 31668 15148 31724
rect 8418 31612 8428 31668
rect 8484 31612 10892 31668
rect 10948 31612 15148 31668
rect 15250 31612 15260 31668
rect 15316 31612 17836 31668
rect 17892 31612 17902 31668
rect 19506 31612 19516 31668
rect 19572 31612 21420 31668
rect 21476 31612 21486 31668
rect 23090 31612 23100 31668
rect 23156 31612 32620 31668
rect 32676 31612 32686 31668
rect 35186 31612 35196 31668
rect 35252 31612 35644 31668
rect 35700 31612 37436 31668
rect 37492 31612 37502 31668
rect 12898 31500 12908 31556
rect 12964 31500 17052 31556
rect 17108 31500 17118 31556
rect 18162 31500 18172 31556
rect 18228 31500 20300 31556
rect 20356 31500 20366 31556
rect 20626 31500 20636 31556
rect 20692 31500 21868 31556
rect 21924 31500 21934 31556
rect 24434 31500 24444 31556
rect 24500 31500 29708 31556
rect 29764 31500 29774 31556
rect 30930 31500 30940 31556
rect 30996 31500 37212 31556
rect 37268 31500 37278 31556
rect 9090 31388 9100 31444
rect 9156 31388 9436 31444
rect 9492 31388 9502 31444
rect 10994 31388 11004 31444
rect 11060 31388 17332 31444
rect 17714 31388 17724 31444
rect 17780 31388 18508 31444
rect 18564 31388 18574 31444
rect 18834 31388 18844 31444
rect 18900 31388 18956 31444
rect 19012 31388 19292 31444
rect 19348 31388 19358 31444
rect 17276 31332 17332 31388
rect 19826 31332 19836 31388
rect 19892 31332 19940 31388
rect 19996 31332 20044 31388
rect 20100 31332 20110 31388
rect 50546 31332 50556 31388
rect 50612 31332 50660 31388
rect 50716 31332 50764 31388
rect 50820 31332 50830 31388
rect 6066 31276 6076 31332
rect 6132 31276 7420 31332
rect 7476 31276 7486 31332
rect 13122 31276 13132 31332
rect 13188 31276 13804 31332
rect 13860 31276 17052 31332
rect 17108 31276 17118 31332
rect 17266 31276 17276 31332
rect 17332 31276 17612 31332
rect 17668 31276 17678 31332
rect 21410 31276 21420 31332
rect 21476 31276 22652 31332
rect 22708 31276 22718 31332
rect 23202 31276 23212 31332
rect 23268 31276 25900 31332
rect 25956 31276 26124 31332
rect 26180 31276 26190 31332
rect 2034 31164 2044 31220
rect 2100 31164 2110 31220
rect 5506 31164 5516 31220
rect 5572 31164 5964 31220
rect 6020 31164 6030 31220
rect 7522 31164 7532 31220
rect 7588 31164 15036 31220
rect 15092 31164 15102 31220
rect 15362 31164 15372 31220
rect 15428 31164 16156 31220
rect 16212 31164 16222 31220
rect 18022 31164 18060 31220
rect 18116 31164 18126 31220
rect 18694 31164 18732 31220
rect 18788 31164 18798 31220
rect 19058 31164 19068 31220
rect 19124 31164 19740 31220
rect 19796 31164 19806 31220
rect 23874 31164 23884 31220
rect 23940 31164 26348 31220
rect 26404 31164 26414 31220
rect 27794 31164 27804 31220
rect 27860 31164 29372 31220
rect 29428 31164 29438 31220
rect 29698 31164 29708 31220
rect 29764 31164 33180 31220
rect 33236 31164 33246 31220
rect 2044 31108 2100 31164
rect 2044 31052 3052 31108
rect 3108 31052 3118 31108
rect 7532 30996 7588 31164
rect 12562 31052 12572 31108
rect 12628 31052 13468 31108
rect 13524 31052 13534 31108
rect 14214 31052 14252 31108
rect 14308 31052 14318 31108
rect 14466 31052 14476 31108
rect 14532 31052 14570 31108
rect 15474 31052 15484 31108
rect 15540 31052 15708 31108
rect 15764 31052 15774 31108
rect 16268 31052 17612 31108
rect 17668 31052 17678 31108
rect 18834 31052 18844 31108
rect 18900 31052 24444 31108
rect 24500 31052 24510 31108
rect 34178 31052 34188 31108
rect 34244 31052 34412 31108
rect 34468 31052 35756 31108
rect 35812 31052 39452 31108
rect 39508 31052 39518 31108
rect 5506 30940 5516 30996
rect 5572 30940 5964 30996
rect 6020 30940 7588 30996
rect 8978 30940 8988 30996
rect 9044 30940 10108 30996
rect 10164 30940 11116 30996
rect 11172 30940 11182 30996
rect 14130 30940 14140 30996
rect 14196 30940 15260 30996
rect 15316 30940 15326 30996
rect 15484 30884 15540 31052
rect 16268 30996 16324 31052
rect 16034 30940 16044 30996
rect 16100 30940 16268 30996
rect 16324 30940 16334 30996
rect 16818 30940 16828 30996
rect 16884 30940 17836 30996
rect 17892 30940 18956 30996
rect 19012 30940 19022 30996
rect 24210 30940 24220 30996
rect 24276 30940 26236 30996
rect 26292 30940 26302 30996
rect 33730 30940 33740 30996
rect 33796 30940 35980 30996
rect 36036 30940 36876 30996
rect 36932 30940 36942 30996
rect 3378 30828 3388 30884
rect 3444 30828 4396 30884
rect 4452 30828 4462 30884
rect 12114 30828 12124 30884
rect 12180 30828 15540 30884
rect 17154 30828 17164 30884
rect 17220 30828 19292 30884
rect 19348 30828 23212 30884
rect 23268 30828 23278 30884
rect 26852 30828 27132 30884
rect 27188 30828 28028 30884
rect 28084 30828 28094 30884
rect 0 30772 800 30800
rect 26852 30772 26908 30828
rect 0 30716 1708 30772
rect 1764 30716 1774 30772
rect 13010 30716 13020 30772
rect 13076 30716 14924 30772
rect 14980 30716 14990 30772
rect 20066 30716 20076 30772
rect 20132 30716 21420 30772
rect 21476 30716 26908 30772
rect 0 30688 800 30716
rect 14130 30604 14140 30660
rect 14196 30604 15036 30660
rect 15092 30604 15102 30660
rect 19282 30604 19292 30660
rect 19348 30604 25676 30660
rect 25732 30604 25742 30660
rect 4466 30548 4476 30604
rect 4532 30548 4580 30604
rect 4636 30548 4684 30604
rect 4740 30548 4750 30604
rect 35186 30548 35196 30604
rect 35252 30548 35300 30604
rect 35356 30548 35404 30604
rect 35460 30548 35470 30604
rect 11414 30492 11452 30548
rect 11508 30492 11518 30548
rect 16034 30492 16044 30548
rect 16100 30492 16268 30548
rect 16324 30492 16334 30548
rect 17938 30492 17948 30548
rect 18004 30492 27692 30548
rect 27748 30492 27758 30548
rect 11218 30380 11228 30436
rect 11284 30380 11564 30436
rect 11620 30380 11630 30436
rect 14578 30380 14588 30436
rect 14644 30380 19964 30436
rect 20020 30380 20030 30436
rect 21410 30380 21420 30436
rect 21476 30380 21756 30436
rect 21812 30380 21822 30436
rect 25862 30380 25900 30436
rect 25956 30380 28364 30436
rect 28420 30380 28700 30436
rect 28756 30380 28766 30436
rect 7970 30268 7980 30324
rect 8036 30268 11900 30324
rect 11956 30268 11966 30324
rect 14354 30268 14364 30324
rect 14420 30268 20972 30324
rect 21028 30268 21038 30324
rect 28018 30268 28028 30324
rect 28084 30268 31500 30324
rect 31556 30268 31566 30324
rect 6636 30156 16156 30212
rect 16212 30156 17724 30212
rect 17780 30156 18732 30212
rect 18788 30156 18798 30212
rect 20738 30156 20748 30212
rect 20804 30156 23548 30212
rect 23604 30156 23614 30212
rect 24546 30156 24556 30212
rect 24612 30156 25228 30212
rect 25284 30156 26796 30212
rect 26852 30156 26862 30212
rect 27570 30156 27580 30212
rect 27636 30156 28028 30212
rect 28084 30156 28094 30212
rect 30930 30156 30940 30212
rect 30996 30156 31948 30212
rect 32004 30156 32014 30212
rect 34962 30156 34972 30212
rect 35028 30156 35644 30212
rect 35700 30156 36988 30212
rect 37044 30156 37054 30212
rect 37202 30156 37212 30212
rect 37268 30156 38108 30212
rect 38164 30156 38174 30212
rect 6636 30100 6692 30156
rect 37212 30100 37268 30156
rect 2034 30044 2044 30100
rect 2100 30044 6188 30100
rect 6244 30044 6254 30100
rect 6626 30044 6636 30100
rect 6692 30044 6702 30100
rect 8642 30044 8652 30100
rect 8708 30044 11788 30100
rect 11844 30044 11854 30100
rect 12114 30044 12124 30100
rect 12180 30044 13692 30100
rect 13748 30044 13758 30100
rect 14886 30044 14924 30100
rect 14980 30044 14990 30100
rect 16482 30044 16492 30100
rect 16548 30044 17276 30100
rect 17332 30044 17342 30100
rect 19954 30044 19964 30100
rect 20020 30044 20300 30100
rect 20356 30044 22540 30100
rect 22596 30044 22606 30100
rect 23202 30044 23212 30100
rect 23268 30044 24108 30100
rect 24164 30044 25116 30100
rect 25172 30044 25182 30100
rect 30482 30044 30492 30100
rect 30548 30044 31052 30100
rect 31108 30044 31118 30100
rect 35970 30044 35980 30100
rect 36036 30044 36540 30100
rect 36596 30044 37268 30100
rect 11732 29988 11788 30044
rect 2370 29932 2380 29988
rect 2436 29932 3164 29988
rect 3220 29932 3230 29988
rect 4162 29932 4172 29988
rect 4228 29932 5068 29988
rect 5124 29932 5134 29988
rect 5730 29932 5740 29988
rect 5796 29932 5852 29988
rect 5908 29932 5918 29988
rect 7746 29932 7756 29988
rect 7812 29932 9996 29988
rect 10052 29932 10062 29988
rect 10434 29932 10444 29988
rect 10500 29932 10892 29988
rect 10948 29932 10958 29988
rect 11106 29932 11116 29988
rect 11172 29932 11564 29988
rect 11620 29932 11630 29988
rect 11732 29932 12684 29988
rect 12740 29932 12750 29988
rect 15138 29932 15148 29988
rect 15204 29932 15242 29988
rect 19628 29932 20076 29988
rect 20132 29932 20142 29988
rect 23538 29932 23548 29988
rect 23604 29932 25340 29988
rect 25396 29932 25406 29988
rect 26002 29932 26012 29988
rect 26068 29932 27748 29988
rect 27906 29932 27916 29988
rect 27972 29932 29260 29988
rect 29316 29932 29326 29988
rect 32834 29932 32844 29988
rect 32900 29932 32910 29988
rect 3714 29820 3724 29876
rect 3780 29820 6412 29876
rect 6468 29820 7868 29876
rect 7924 29820 7934 29876
rect 9650 29820 9660 29876
rect 9716 29820 10668 29876
rect 10724 29820 13580 29876
rect 13636 29820 13646 29876
rect 18162 29820 18172 29876
rect 18228 29820 18396 29876
rect 18452 29820 18956 29876
rect 19012 29820 19022 29876
rect 1138 29708 1148 29764
rect 1204 29708 7532 29764
rect 7588 29708 7598 29764
rect 11218 29708 11228 29764
rect 11284 29708 11900 29764
rect 11956 29708 11966 29764
rect 12450 29708 12460 29764
rect 12516 29708 13356 29764
rect 13412 29708 19068 29764
rect 19124 29708 19134 29764
rect 19628 29652 19684 29932
rect 27692 29876 27748 29932
rect 32844 29876 32900 29932
rect 22642 29820 22652 29876
rect 22708 29820 23436 29876
rect 23492 29820 27188 29876
rect 27692 29820 32900 29876
rect 19826 29764 19836 29820
rect 19892 29764 19940 29820
rect 19996 29764 20044 29820
rect 20100 29764 20110 29820
rect 21186 29708 21196 29764
rect 21252 29708 23884 29764
rect 23940 29708 24332 29764
rect 24388 29708 25956 29764
rect 19628 29596 19740 29652
rect 19796 29596 19806 29652
rect 20066 29596 20076 29652
rect 20132 29596 21308 29652
rect 21364 29596 21374 29652
rect 21970 29596 21980 29652
rect 22036 29596 24108 29652
rect 24164 29596 25564 29652
rect 25620 29596 25630 29652
rect 19628 29540 19684 29596
rect 5618 29484 5628 29540
rect 5684 29484 7420 29540
rect 7476 29484 7486 29540
rect 11778 29484 11788 29540
rect 11844 29484 19684 29540
rect 20402 29484 20412 29540
rect 20468 29484 21084 29540
rect 21140 29484 22428 29540
rect 22484 29484 22494 29540
rect 4610 29372 4620 29428
rect 4676 29372 5740 29428
rect 5796 29372 5806 29428
rect 9650 29372 9660 29428
rect 9716 29372 10668 29428
rect 10724 29372 10734 29428
rect 10994 29372 11004 29428
rect 11060 29372 11900 29428
rect 11956 29372 11966 29428
rect 12114 29372 12124 29428
rect 12180 29372 14812 29428
rect 14868 29372 14878 29428
rect 18722 29372 18732 29428
rect 18788 29372 20972 29428
rect 21028 29372 21038 29428
rect 21522 29372 21532 29428
rect 21588 29372 21980 29428
rect 22036 29372 23100 29428
rect 23156 29372 23166 29428
rect 12124 29316 12180 29372
rect 25900 29316 25956 29708
rect 27132 29652 27188 29820
rect 50546 29764 50556 29820
rect 50612 29764 50660 29820
rect 50716 29764 50764 29820
rect 50820 29764 50830 29820
rect 27122 29596 27132 29652
rect 27188 29596 27692 29652
rect 27748 29596 30268 29652
rect 30324 29596 30334 29652
rect 28354 29372 28364 29428
rect 28420 29372 28924 29428
rect 28980 29372 29708 29428
rect 29764 29372 29774 29428
rect 2818 29260 2828 29316
rect 2884 29260 3164 29316
rect 3220 29260 3230 29316
rect 5058 29260 5068 29316
rect 5124 29260 8540 29316
rect 8596 29260 12180 29316
rect 12646 29260 12684 29316
rect 12740 29260 12750 29316
rect 13682 29260 13692 29316
rect 13748 29260 24444 29316
rect 24500 29260 25676 29316
rect 25732 29260 25742 29316
rect 25900 29260 27356 29316
rect 27412 29260 27422 29316
rect 27794 29260 27804 29316
rect 27860 29260 29596 29316
rect 29652 29260 29662 29316
rect 14242 29148 14252 29204
rect 14308 29148 14318 29204
rect 19058 29148 19068 29204
rect 19124 29148 20076 29204
rect 20132 29148 20142 29204
rect 26002 29148 26012 29204
rect 26068 29148 26908 29204
rect 26964 29148 30492 29204
rect 30548 29148 30558 29204
rect 14252 29092 14308 29148
rect 14252 29036 20188 29092
rect 20244 29036 20254 29092
rect 0 28980 800 29008
rect 4466 28980 4476 29036
rect 4532 28980 4580 29036
rect 4636 28980 4684 29036
rect 4740 28980 4750 29036
rect 35186 28980 35196 29036
rect 35252 28980 35300 29036
rect 35356 28980 35404 29036
rect 35460 28980 35470 29036
rect 0 28924 2380 28980
rect 2436 28924 2446 28980
rect 18610 28924 18620 28980
rect 18676 28924 19964 28980
rect 20020 28924 20030 28980
rect 0 28896 800 28924
rect 9090 28812 9100 28868
rect 9156 28812 11340 28868
rect 11396 28812 12236 28868
rect 12292 28812 18732 28868
rect 18788 28812 19236 28868
rect 19394 28812 19404 28868
rect 19460 28812 26684 28868
rect 26740 28812 27244 28868
rect 27300 28812 27310 28868
rect 19180 28756 19236 28812
rect 12674 28700 12684 28756
rect 12740 28700 13356 28756
rect 13412 28700 13422 28756
rect 14326 28700 14364 28756
rect 14420 28700 15260 28756
rect 15316 28700 15326 28756
rect 16706 28700 16716 28756
rect 16772 28700 17500 28756
rect 17556 28700 17566 28756
rect 19170 28700 19180 28756
rect 19236 28700 26348 28756
rect 26404 28700 26414 28756
rect 27346 28700 27356 28756
rect 27412 28700 28252 28756
rect 28308 28700 28318 28756
rect 28466 28700 28476 28756
rect 28532 28700 29148 28756
rect 29204 28700 29214 28756
rect 2370 28588 2380 28644
rect 2436 28588 2940 28644
rect 2996 28588 3948 28644
rect 4004 28588 5740 28644
rect 5796 28588 5806 28644
rect 8614 28588 8652 28644
rect 8708 28588 8718 28644
rect 8866 28588 8876 28644
rect 8932 28588 10556 28644
rect 10612 28588 18844 28644
rect 18900 28588 18910 28644
rect 23426 28588 23436 28644
rect 23492 28588 25116 28644
rect 25172 28588 26012 28644
rect 26068 28588 26078 28644
rect 18844 28532 18900 28588
rect 2034 28476 2044 28532
rect 2100 28476 3276 28532
rect 3332 28476 3342 28532
rect 5282 28476 5292 28532
rect 5348 28476 7756 28532
rect 7812 28476 7822 28532
rect 8764 28476 12572 28532
rect 12628 28476 12638 28532
rect 13234 28476 13244 28532
rect 13300 28476 14700 28532
rect 14756 28476 14766 28532
rect 14914 28476 14924 28532
rect 14980 28476 16716 28532
rect 16772 28476 16782 28532
rect 18844 28476 21532 28532
rect 21588 28476 21598 28532
rect 22866 28476 22876 28532
rect 22932 28476 24220 28532
rect 24276 28476 24286 28532
rect 8764 28420 8820 28476
rect 1810 28364 1820 28420
rect 1876 28364 2492 28420
rect 2548 28364 2558 28420
rect 2706 28364 2716 28420
rect 2772 28364 3500 28420
rect 3556 28364 3566 28420
rect 5954 28364 5964 28420
rect 6020 28364 8764 28420
rect 8820 28364 8830 28420
rect 10882 28364 10892 28420
rect 10948 28364 15372 28420
rect 15428 28364 15438 28420
rect 16034 28364 16044 28420
rect 16100 28364 18172 28420
rect 18228 28364 18238 28420
rect 19618 28364 19628 28420
rect 19684 28364 20188 28420
rect 20244 28364 20254 28420
rect 24322 28364 24332 28420
rect 24388 28364 28700 28420
rect 28756 28364 29260 28420
rect 29316 28364 29326 28420
rect 1474 28252 1484 28308
rect 1540 28252 4844 28308
rect 4900 28252 5852 28308
rect 5908 28252 5918 28308
rect 8530 28252 8540 28308
rect 8596 28252 8876 28308
rect 8932 28252 8942 28308
rect 19826 28196 19836 28252
rect 19892 28196 19940 28252
rect 19996 28196 20044 28252
rect 20100 28196 20110 28252
rect 50546 28196 50556 28252
rect 50612 28196 50660 28252
rect 50716 28196 50764 28252
rect 50820 28196 50830 28252
rect 7868 28140 17556 28196
rect 3938 28028 3948 28084
rect 4004 28028 5292 28084
rect 5348 28028 5358 28084
rect 7868 27972 7924 28140
rect 8642 28028 8652 28084
rect 8708 28028 9772 28084
rect 9828 28028 9838 28084
rect 10546 28028 10556 28084
rect 10612 28028 11116 28084
rect 11172 28028 11564 28084
rect 11620 28028 12236 28084
rect 12292 28028 13972 28084
rect 14130 28028 14140 28084
rect 14196 28028 15036 28084
rect 15092 28028 15102 28084
rect 15586 28028 15596 28084
rect 15652 28028 15662 28084
rect 4946 27916 4956 27972
rect 5012 27916 6412 27972
rect 6468 27916 7924 27972
rect 13916 27860 13972 28028
rect 15596 27972 15652 28028
rect 15138 27916 15148 27972
rect 15204 27916 16716 27972
rect 16772 27916 16782 27972
rect 17500 27860 17556 28140
rect 23492 28140 30828 28196
rect 30884 28140 30894 28196
rect 23492 27972 23548 28140
rect 24658 28028 24668 28084
rect 24724 28028 25340 28084
rect 25396 28028 25406 28084
rect 29698 28028 29708 28084
rect 29764 28028 30604 28084
rect 30660 28028 35756 28084
rect 35812 28028 35822 28084
rect 19282 27916 19292 27972
rect 19348 27916 20524 27972
rect 20580 27916 20590 27972
rect 21634 27916 21644 27972
rect 21700 27916 23548 27972
rect 27020 27916 27356 27972
rect 27412 27916 27422 27972
rect 27020 27860 27076 27916
rect 5394 27804 5404 27860
rect 5460 27804 7084 27860
rect 7140 27804 7150 27860
rect 7746 27804 7756 27860
rect 7812 27804 10108 27860
rect 10164 27804 10780 27860
rect 10836 27804 10846 27860
rect 12086 27804 12124 27860
rect 12180 27804 12190 27860
rect 12674 27804 12684 27860
rect 12740 27804 13244 27860
rect 13300 27804 13310 27860
rect 13916 27804 14532 27860
rect 15026 27804 15036 27860
rect 15092 27804 15484 27860
rect 15540 27804 15550 27860
rect 17490 27804 17500 27860
rect 17556 27804 17836 27860
rect 17892 27804 18508 27860
rect 18564 27804 19404 27860
rect 19460 27804 19470 27860
rect 19954 27804 19964 27860
rect 20020 27804 25228 27860
rect 25284 27804 26684 27860
rect 26740 27804 27076 27860
rect 27906 27804 27916 27860
rect 27972 27804 30044 27860
rect 30100 27804 30110 27860
rect 14476 27748 14532 27804
rect 1698 27692 1708 27748
rect 1764 27692 2492 27748
rect 2548 27692 2558 27748
rect 5506 27692 5516 27748
rect 5572 27692 5964 27748
rect 6020 27692 6030 27748
rect 8614 27692 8652 27748
rect 8708 27692 8718 27748
rect 8978 27692 8988 27748
rect 9044 27692 9996 27748
rect 10052 27692 14252 27748
rect 14308 27692 14318 27748
rect 14476 27692 22484 27748
rect 22642 27692 22652 27748
rect 22708 27692 23548 27748
rect 23604 27692 23614 27748
rect 26450 27692 26460 27748
rect 26516 27692 28140 27748
rect 28196 27692 28206 27748
rect 22428 27636 22484 27692
rect 4274 27580 4284 27636
rect 4340 27580 15148 27636
rect 15810 27580 15820 27636
rect 15876 27580 16716 27636
rect 16772 27580 16782 27636
rect 18386 27580 18396 27636
rect 18452 27580 19068 27636
rect 19124 27580 19134 27636
rect 22428 27580 24668 27636
rect 24724 27580 25452 27636
rect 25508 27580 25518 27636
rect 7970 27468 7980 27524
rect 8036 27468 8540 27524
rect 8596 27468 14252 27524
rect 14308 27468 14318 27524
rect 4466 27412 4476 27468
rect 4532 27412 4580 27468
rect 4636 27412 4684 27468
rect 4740 27412 4750 27468
rect 15092 27412 15148 27580
rect 16258 27468 16268 27524
rect 16324 27468 20188 27524
rect 20244 27468 20254 27524
rect 35186 27412 35196 27468
rect 35252 27412 35300 27468
rect 35356 27412 35404 27468
rect 35460 27412 35470 27468
rect 15092 27356 18060 27412
rect 18116 27356 18126 27412
rect 12338 27244 12348 27300
rect 12404 27244 14476 27300
rect 14532 27244 16268 27300
rect 16324 27244 16334 27300
rect 17154 27244 17164 27300
rect 17220 27244 28588 27300
rect 28644 27244 29148 27300
rect 29204 27244 29214 27300
rect 0 27188 800 27216
rect 0 27132 1708 27188
rect 1764 27132 1774 27188
rect 6738 27132 6748 27188
rect 6804 27132 9212 27188
rect 9268 27132 9278 27188
rect 14802 27132 14812 27188
rect 14868 27132 15708 27188
rect 15764 27132 15774 27188
rect 17938 27132 17948 27188
rect 18004 27132 18732 27188
rect 18788 27132 18798 27188
rect 21970 27132 21980 27188
rect 22036 27132 23772 27188
rect 23828 27132 24220 27188
rect 24276 27132 24286 27188
rect 0 27104 800 27132
rect 21980 27076 22036 27132
rect 5926 27020 5964 27076
rect 6020 27020 6030 27076
rect 9090 27020 9100 27076
rect 9156 27020 10556 27076
rect 10612 27020 10622 27076
rect 11666 27020 11676 27076
rect 11732 27020 12236 27076
rect 12292 27020 13580 27076
rect 13636 27020 17612 27076
rect 17668 27020 17678 27076
rect 18162 27020 18172 27076
rect 18228 27020 22036 27076
rect 1138 26908 1148 26964
rect 1204 26908 3388 26964
rect 3444 26908 3454 26964
rect 5702 26908 5740 26964
rect 5796 26908 5806 26964
rect 9762 26908 9772 26964
rect 9828 26908 10108 26964
rect 10164 26908 13412 26964
rect 15138 26908 15148 26964
rect 15204 26908 18284 26964
rect 18340 26908 21420 26964
rect 21476 26908 21486 26964
rect 13356 26852 13412 26908
rect 9314 26796 9324 26852
rect 9380 26796 9548 26852
rect 9604 26796 9614 26852
rect 11750 26796 11788 26852
rect 11844 26796 11854 26852
rect 13356 26796 15036 26852
rect 15092 26796 15102 26852
rect 15698 26796 15708 26852
rect 15764 26796 16380 26852
rect 16436 26796 16446 26852
rect 16594 26796 16604 26852
rect 16660 26796 16940 26852
rect 16996 26796 17006 26852
rect 17602 26796 17612 26852
rect 17668 26796 20300 26852
rect 20356 26796 20366 26852
rect 12674 26684 12684 26740
rect 12740 26684 15596 26740
rect 15652 26684 15662 26740
rect 15820 26684 18340 26740
rect 11414 26572 11452 26628
rect 11508 26572 12012 26628
rect 12068 26572 13692 26628
rect 13748 26572 15260 26628
rect 15316 26572 15326 26628
rect 15820 26516 15876 26684
rect 6066 26460 6076 26516
rect 6132 26460 9660 26516
rect 9716 26460 9726 26516
rect 9874 26460 9884 26516
rect 9940 26460 10556 26516
rect 10612 26460 10622 26516
rect 12786 26460 12796 26516
rect 12852 26460 13244 26516
rect 13300 26460 13310 26516
rect 15026 26460 15036 26516
rect 15092 26460 15372 26516
rect 15428 26460 15876 26516
rect 15932 26572 17948 26628
rect 18004 26572 18014 26628
rect 15932 26404 15988 26572
rect 18284 26516 18340 26684
rect 19826 26628 19836 26684
rect 19892 26628 19940 26684
rect 19996 26628 20044 26684
rect 20100 26628 20110 26684
rect 50546 26628 50556 26684
rect 50612 26628 50660 26684
rect 50716 26628 50764 26684
rect 50820 26628 50830 26684
rect 20178 26572 20188 26628
rect 20244 26572 27804 26628
rect 27860 26572 28252 26628
rect 28308 26572 28318 26628
rect 18284 26460 21084 26516
rect 21140 26460 21150 26516
rect 7858 26348 7868 26404
rect 7924 26348 8428 26404
rect 10210 26348 10220 26404
rect 10276 26348 11004 26404
rect 11060 26348 11070 26404
rect 13906 26348 13916 26404
rect 13972 26348 15988 26404
rect 16146 26348 16156 26404
rect 16212 26348 17612 26404
rect 17668 26348 18508 26404
rect 18564 26348 25508 26404
rect 5954 26236 5964 26292
rect 6020 26236 7644 26292
rect 7700 26236 7710 26292
rect 8372 26068 8428 26348
rect 15708 26292 15764 26348
rect 25452 26292 25508 26348
rect 9650 26236 9660 26292
rect 9716 26236 11900 26292
rect 11956 26236 13580 26292
rect 13636 26236 13646 26292
rect 15698 26236 15708 26292
rect 15764 26236 15774 26292
rect 16034 26236 16044 26292
rect 16100 26236 17948 26292
rect 18004 26236 18014 26292
rect 21634 26236 21644 26292
rect 21700 26236 22092 26292
rect 22148 26236 23100 26292
rect 23156 26236 23166 26292
rect 25442 26236 25452 26292
rect 25508 26236 26796 26292
rect 26852 26236 26862 26292
rect 10546 26124 10556 26180
rect 10612 26124 16380 26180
rect 16436 26124 16940 26180
rect 16996 26124 17388 26180
rect 17444 26124 17454 26180
rect 19170 26124 19180 26180
rect 19236 26124 19852 26180
rect 19908 26124 19918 26180
rect 20738 26124 20748 26180
rect 20804 26124 25564 26180
rect 25620 26124 25630 26180
rect 19180 26068 19236 26124
rect 8372 26012 19236 26068
rect 10994 25900 11004 25956
rect 11060 25900 15932 25956
rect 15988 25900 15998 25956
rect 4466 25844 4476 25900
rect 4532 25844 4580 25900
rect 4636 25844 4684 25900
rect 4740 25844 4750 25900
rect 35186 25844 35196 25900
rect 35252 25844 35300 25900
rect 35356 25844 35404 25900
rect 35460 25844 35470 25900
rect 14130 25788 14140 25844
rect 14196 25788 14476 25844
rect 14532 25788 14924 25844
rect 14980 25788 17612 25844
rect 17668 25788 19964 25844
rect 20020 25788 20030 25844
rect 20412 25788 23324 25844
rect 23380 25788 24444 25844
rect 24500 25788 24510 25844
rect 20412 25732 20468 25788
rect 6850 25676 6860 25732
rect 6916 25676 7308 25732
rect 7364 25676 7374 25732
rect 9538 25676 9548 25732
rect 9604 25676 14756 25732
rect 15810 25676 15820 25732
rect 15876 25676 16268 25732
rect 16324 25676 20468 25732
rect 22754 25676 22764 25732
rect 22820 25676 23548 25732
rect 23604 25676 23614 25732
rect 7074 25564 7084 25620
rect 7140 25564 7756 25620
rect 7812 25564 9660 25620
rect 9716 25564 9726 25620
rect 14700 25508 14756 25676
rect 16044 25564 16716 25620
rect 16772 25564 16782 25620
rect 19730 25564 19740 25620
rect 19796 25564 20300 25620
rect 20356 25564 25340 25620
rect 25396 25564 27132 25620
rect 27188 25564 33628 25620
rect 33684 25564 33694 25620
rect 16044 25508 16100 25564
rect 7522 25452 7532 25508
rect 7588 25452 10220 25508
rect 10276 25452 10286 25508
rect 10994 25452 11004 25508
rect 11060 25452 11900 25508
rect 11956 25452 11966 25508
rect 14690 25452 14700 25508
rect 14756 25452 16044 25508
rect 16100 25452 16110 25508
rect 16818 25452 16828 25508
rect 16884 25452 18844 25508
rect 18900 25452 19404 25508
rect 19460 25452 19470 25508
rect 19842 25452 19852 25508
rect 19908 25452 23660 25508
rect 23716 25452 23726 25508
rect 0 25396 800 25424
rect 0 25340 1708 25396
rect 1764 25340 2492 25396
rect 2548 25340 2558 25396
rect 9538 25340 9548 25396
rect 9604 25340 10444 25396
rect 10500 25340 10510 25396
rect 10770 25340 10780 25396
rect 10836 25340 12572 25396
rect 12628 25340 12638 25396
rect 15586 25340 15596 25396
rect 15652 25340 16156 25396
rect 16212 25340 20188 25396
rect 20244 25340 20254 25396
rect 22642 25340 22652 25396
rect 22708 25340 23548 25396
rect 23604 25340 23614 25396
rect 0 25312 800 25340
rect 7858 25228 7868 25284
rect 7924 25228 8316 25284
rect 8372 25228 11676 25284
rect 11732 25228 11742 25284
rect 12450 25228 12460 25284
rect 12516 25228 13468 25284
rect 13524 25228 13916 25284
rect 13972 25228 13982 25284
rect 17714 25228 17724 25284
rect 17780 25228 18620 25284
rect 18676 25228 18686 25284
rect 19058 25228 19068 25284
rect 19124 25228 20076 25284
rect 20132 25228 21532 25284
rect 21588 25228 22540 25284
rect 22596 25228 22606 25284
rect 27794 25228 27804 25284
rect 27860 25228 29260 25284
rect 29316 25228 36428 25284
rect 36484 25228 36494 25284
rect 14018 25116 14028 25172
rect 14084 25116 17388 25172
rect 17444 25116 17454 25172
rect 19068 25060 19124 25228
rect 23090 25116 23100 25172
rect 23156 25116 24444 25172
rect 24500 25116 24510 25172
rect 19826 25060 19836 25116
rect 19892 25060 19940 25116
rect 19996 25060 20044 25116
rect 20100 25060 20110 25116
rect 50546 25060 50556 25116
rect 50612 25060 50660 25116
rect 50716 25060 50764 25116
rect 50820 25060 50830 25116
rect 1474 25004 1484 25060
rect 1540 25004 4732 25060
rect 4788 25004 4798 25060
rect 8194 25004 8204 25060
rect 8260 25004 19124 25060
rect 11666 24892 11676 24948
rect 11732 24892 12348 24948
rect 12404 24892 12414 24948
rect 17266 24892 17276 24948
rect 17332 24892 22372 24948
rect 25778 24892 25788 24948
rect 25844 24892 26236 24948
rect 26292 24892 32060 24948
rect 32116 24892 32126 24948
rect 22316 24836 22372 24892
rect 13346 24780 13356 24836
rect 13412 24780 14252 24836
rect 14308 24780 22092 24836
rect 22148 24780 22158 24836
rect 22316 24780 30492 24836
rect 30548 24780 30558 24836
rect 11666 24668 11676 24724
rect 11732 24668 16492 24724
rect 16548 24668 16558 24724
rect 16706 24668 16716 24724
rect 16772 24668 17836 24724
rect 17892 24668 19964 24724
rect 20020 24668 20030 24724
rect 22194 24668 22204 24724
rect 22260 24668 24220 24724
rect 24276 24668 25004 24724
rect 25060 24668 25070 24724
rect 16492 24612 16548 24668
rect 16492 24556 16828 24612
rect 16884 24556 16894 24612
rect 18470 24556 18508 24612
rect 18564 24556 18574 24612
rect 19058 24556 19068 24612
rect 19124 24556 24108 24612
rect 24164 24556 25228 24612
rect 25284 24556 25294 24612
rect 4466 24276 4476 24332
rect 4532 24276 4580 24332
rect 4636 24276 4684 24332
rect 4740 24276 4750 24332
rect 35186 24276 35196 24332
rect 35252 24276 35300 24332
rect 35356 24276 35404 24332
rect 35460 24276 35470 24332
rect 12898 24220 12908 24276
rect 12964 24220 14700 24276
rect 14756 24220 23772 24276
rect 23828 24220 24332 24276
rect 24388 24220 24398 24276
rect 11330 24108 11340 24164
rect 11396 24108 15708 24164
rect 15764 24108 15774 24164
rect 19516 24108 22316 24164
rect 22372 24108 22382 24164
rect 19516 24052 19572 24108
rect 9874 23996 9884 24052
rect 9940 23996 15148 24052
rect 15204 23996 19572 24052
rect 19730 23996 19740 24052
rect 19796 23996 20524 24052
rect 20580 23996 20590 24052
rect 24434 23996 24444 24052
rect 24500 23996 25788 24052
rect 25844 23996 25854 24052
rect 15446 23884 15484 23940
rect 15540 23884 15550 23940
rect 20178 23884 20188 23940
rect 20244 23884 21084 23940
rect 21140 23884 21150 23940
rect 24770 23884 24780 23940
rect 24836 23884 25452 23940
rect 25508 23884 25518 23940
rect 2034 23772 2044 23828
rect 2100 23772 3164 23828
rect 3220 23772 3230 23828
rect 15810 23772 15820 23828
rect 15876 23772 18172 23828
rect 18228 23772 21532 23828
rect 21588 23772 21598 23828
rect 0 23604 800 23632
rect 0 23548 1708 23604
rect 1764 23548 2492 23604
rect 2548 23548 2558 23604
rect 21074 23548 21084 23604
rect 21140 23548 21868 23604
rect 21924 23548 21934 23604
rect 0 23520 800 23548
rect 19826 23492 19836 23548
rect 19892 23492 19940 23548
rect 19996 23492 20044 23548
rect 20100 23492 20110 23548
rect 50546 23492 50556 23548
rect 50612 23492 50660 23548
rect 50716 23492 50764 23548
rect 50820 23492 50830 23548
rect 1026 23436 1036 23492
rect 1092 23436 2380 23492
rect 2436 23436 2446 23492
rect 20188 23436 23996 23492
rect 24052 23436 24062 23492
rect 20188 23380 20244 23436
rect 10322 23324 10332 23380
rect 10388 23324 20244 23380
rect 22194 23324 22204 23380
rect 22260 23324 22988 23380
rect 23044 23324 23054 23380
rect 5842 23212 5852 23268
rect 5908 23212 8428 23268
rect 15810 23212 15820 23268
rect 15876 23212 21308 23268
rect 21364 23212 21374 23268
rect 8372 23156 8428 23212
rect 8372 23100 27020 23156
rect 27076 23100 27086 23156
rect 16146 22876 16156 22932
rect 16212 22876 17612 22932
rect 17668 22876 27916 22932
rect 27972 22876 27982 22932
rect 4466 22708 4476 22764
rect 4532 22708 4580 22764
rect 4636 22708 4684 22764
rect 4740 22708 4750 22764
rect 35186 22708 35196 22764
rect 35252 22708 35300 22764
rect 35356 22708 35404 22764
rect 35460 22708 35470 22764
rect 15138 22652 15148 22708
rect 15204 22652 27804 22708
rect 27860 22652 27870 22708
rect 19826 21924 19836 21980
rect 19892 21924 19940 21980
rect 19996 21924 20044 21980
rect 20100 21924 20110 21980
rect 50546 21924 50556 21980
rect 50612 21924 50660 21980
rect 50716 21924 50764 21980
rect 50820 21924 50830 21980
rect 0 21812 800 21840
rect 0 21756 1708 21812
rect 1764 21756 2492 21812
rect 2548 21756 2558 21812
rect 7970 21756 7980 21812
rect 8036 21756 23100 21812
rect 23156 21756 23166 21812
rect 0 21728 800 21756
rect 12674 21644 12684 21700
rect 12740 21644 27804 21700
rect 27860 21644 27870 21700
rect 4466 21140 4476 21196
rect 4532 21140 4580 21196
rect 4636 21140 4684 21196
rect 4740 21140 4750 21196
rect 35186 21140 35196 21196
rect 35252 21140 35300 21196
rect 35356 21140 35404 21196
rect 35460 21140 35470 21196
rect 19826 20356 19836 20412
rect 19892 20356 19940 20412
rect 19996 20356 20044 20412
rect 20100 20356 20110 20412
rect 50546 20356 50556 20412
rect 50612 20356 50660 20412
rect 50716 20356 50764 20412
rect 50820 20356 50830 20412
rect 0 20020 800 20048
rect 0 19964 1708 20020
rect 1764 19964 2492 20020
rect 2548 19964 2558 20020
rect 0 19936 800 19964
rect 4466 19572 4476 19628
rect 4532 19572 4580 19628
rect 4636 19572 4684 19628
rect 4740 19572 4750 19628
rect 35186 19572 35196 19628
rect 35252 19572 35300 19628
rect 35356 19572 35404 19628
rect 35460 19572 35470 19628
rect 19826 18788 19836 18844
rect 19892 18788 19940 18844
rect 19996 18788 20044 18844
rect 20100 18788 20110 18844
rect 50546 18788 50556 18844
rect 50612 18788 50660 18844
rect 50716 18788 50764 18844
rect 50820 18788 50830 18844
rect 0 18228 800 18256
rect 0 18172 1708 18228
rect 1764 18172 2492 18228
rect 2548 18172 2558 18228
rect 0 18144 800 18172
rect 4466 18004 4476 18060
rect 4532 18004 4580 18060
rect 4636 18004 4684 18060
rect 4740 18004 4750 18060
rect 35186 18004 35196 18060
rect 35252 18004 35300 18060
rect 35356 18004 35404 18060
rect 35460 18004 35470 18060
rect 19826 17220 19836 17276
rect 19892 17220 19940 17276
rect 19996 17220 20044 17276
rect 20100 17220 20110 17276
rect 50546 17220 50556 17276
rect 50612 17220 50660 17276
rect 50716 17220 50764 17276
rect 50820 17220 50830 17276
rect 0 16436 800 16464
rect 4466 16436 4476 16492
rect 4532 16436 4580 16492
rect 4636 16436 4684 16492
rect 4740 16436 4750 16492
rect 35186 16436 35196 16492
rect 35252 16436 35300 16492
rect 35356 16436 35404 16492
rect 35460 16436 35470 16492
rect 0 16380 1708 16436
rect 1764 16380 2492 16436
rect 2548 16380 2558 16436
rect 0 16352 800 16380
rect 19826 15652 19836 15708
rect 19892 15652 19940 15708
rect 19996 15652 20044 15708
rect 20100 15652 20110 15708
rect 50546 15652 50556 15708
rect 50612 15652 50660 15708
rect 50716 15652 50764 15708
rect 50820 15652 50830 15708
rect 1138 15148 1148 15204
rect 1204 15148 1820 15204
rect 1876 15148 1886 15204
rect 4466 14868 4476 14924
rect 4532 14868 4580 14924
rect 4636 14868 4684 14924
rect 4740 14868 4750 14924
rect 35186 14868 35196 14924
rect 35252 14868 35300 14924
rect 35356 14868 35404 14924
rect 35460 14868 35470 14924
rect 0 14644 800 14672
rect 0 14588 1708 14644
rect 1764 14588 2492 14644
rect 2548 14588 2558 14644
rect 0 14560 800 14588
rect 19826 14084 19836 14140
rect 19892 14084 19940 14140
rect 19996 14084 20044 14140
rect 20100 14084 20110 14140
rect 50546 14084 50556 14140
rect 50612 14084 50660 14140
rect 50716 14084 50764 14140
rect 50820 14084 50830 14140
rect 2034 13356 2044 13412
rect 2100 13356 3836 13412
rect 3892 13356 3902 13412
rect 4466 13300 4476 13356
rect 4532 13300 4580 13356
rect 4636 13300 4684 13356
rect 4740 13300 4750 13356
rect 35186 13300 35196 13356
rect 35252 13300 35300 13356
rect 35356 13300 35404 13356
rect 35460 13300 35470 13356
rect 0 12852 800 12880
rect 0 12796 1708 12852
rect 1764 12796 2492 12852
rect 2548 12796 2558 12852
rect 0 12768 800 12796
rect 19826 12516 19836 12572
rect 19892 12516 19940 12572
rect 19996 12516 20044 12572
rect 20100 12516 20110 12572
rect 50546 12516 50556 12572
rect 50612 12516 50660 12572
rect 50716 12516 50764 12572
rect 50820 12516 50830 12572
rect 4466 11732 4476 11788
rect 4532 11732 4580 11788
rect 4636 11732 4684 11788
rect 4740 11732 4750 11788
rect 35186 11732 35196 11788
rect 35252 11732 35300 11788
rect 35356 11732 35404 11788
rect 35460 11732 35470 11788
rect 2034 11228 2044 11284
rect 2100 11228 6300 11284
rect 6356 11228 6366 11284
rect 0 11060 800 11088
rect 0 11004 1708 11060
rect 1764 11004 2492 11060
rect 2548 11004 2558 11060
rect 0 10976 800 11004
rect 19826 10948 19836 11004
rect 19892 10948 19940 11004
rect 19996 10948 20044 11004
rect 20100 10948 20110 11004
rect 50546 10948 50556 11004
rect 50612 10948 50660 11004
rect 50716 10948 50764 11004
rect 50820 10948 50830 11004
rect 4466 10164 4476 10220
rect 4532 10164 4580 10220
rect 4636 10164 4684 10220
rect 4740 10164 4750 10220
rect 35186 10164 35196 10220
rect 35252 10164 35300 10220
rect 35356 10164 35404 10220
rect 35460 10164 35470 10220
rect 2370 9996 2380 10052
rect 2436 9996 6524 10052
rect 6580 9996 6590 10052
rect 19826 9380 19836 9436
rect 19892 9380 19940 9436
rect 19996 9380 20044 9436
rect 20100 9380 20110 9436
rect 50546 9380 50556 9436
rect 50612 9380 50660 9436
rect 50716 9380 50764 9436
rect 50820 9380 50830 9436
rect 0 9268 800 9296
rect 0 9212 1708 9268
rect 1764 9212 2492 9268
rect 2548 9212 2558 9268
rect 0 9184 800 9212
rect 4466 8596 4476 8652
rect 4532 8596 4580 8652
rect 4636 8596 4684 8652
rect 4740 8596 4750 8652
rect 35186 8596 35196 8652
rect 35252 8596 35300 8652
rect 35356 8596 35404 8652
rect 35460 8596 35470 8652
rect 1698 7980 1708 8036
rect 1764 7980 2492 8036
rect 2548 7980 2558 8036
rect 19826 7812 19836 7868
rect 19892 7812 19940 7868
rect 19996 7812 20044 7868
rect 20100 7812 20110 7868
rect 50546 7812 50556 7868
rect 50612 7812 50660 7868
rect 50716 7812 50764 7868
rect 50820 7812 50830 7868
rect 0 7476 800 7504
rect 0 7420 1708 7476
rect 1764 7420 1774 7476
rect 0 7392 800 7420
rect 4466 7028 4476 7084
rect 4532 7028 4580 7084
rect 4636 7028 4684 7084
rect 4740 7028 4750 7084
rect 35186 7028 35196 7084
rect 35252 7028 35300 7084
rect 35356 7028 35404 7084
rect 35460 7028 35470 7084
rect 19826 6244 19836 6300
rect 19892 6244 19940 6300
rect 19996 6244 20044 6300
rect 20100 6244 20110 6300
rect 50546 6244 50556 6300
rect 50612 6244 50660 6300
rect 50716 6244 50764 6300
rect 50820 6244 50830 6300
rect 1250 5852 1260 5908
rect 1316 5852 2156 5908
rect 2212 5852 2222 5908
rect 0 5684 800 5712
rect 0 5628 1708 5684
rect 1764 5628 1774 5684
rect 0 5600 800 5628
rect 4466 5460 4476 5516
rect 4532 5460 4580 5516
rect 4636 5460 4684 5516
rect 4740 5460 4750 5516
rect 35186 5460 35196 5516
rect 35252 5460 35300 5516
rect 35356 5460 35404 5516
rect 35460 5460 35470 5516
rect 19826 4676 19836 4732
rect 19892 4676 19940 4732
rect 19996 4676 20044 4732
rect 20100 4676 20110 4732
rect 50546 4676 50556 4732
rect 50612 4676 50660 4732
rect 50716 4676 50764 4732
rect 50820 4676 50830 4732
rect 2034 4508 2044 4564
rect 2100 4508 8204 4564
rect 8260 4508 8270 4564
rect 0 3892 800 3920
rect 4466 3892 4476 3948
rect 4532 3892 4580 3948
rect 4636 3892 4684 3948
rect 4740 3892 4750 3948
rect 35186 3892 35196 3948
rect 35252 3892 35300 3948
rect 35356 3892 35404 3948
rect 35460 3892 35470 3948
rect 0 3836 1708 3892
rect 1764 3836 2492 3892
rect 2548 3836 2558 3892
rect 0 3808 800 3836
rect 1698 3276 1708 3332
rect 1764 3276 2716 3332
rect 2772 3276 2782 3332
rect 19826 3108 19836 3164
rect 19892 3108 19940 3164
rect 19996 3108 20044 3164
rect 20100 3108 20110 3164
rect 50546 3108 50556 3164
rect 50612 3108 50660 3164
rect 50716 3108 50764 3164
rect 50820 3108 50830 3164
rect 0 2100 800 2128
rect 0 2044 1708 2100
rect 1764 2044 1774 2100
rect 0 2016 800 2044
<< via3 >>
rect 19836 56420 19892 56476
rect 19940 56420 19996 56476
rect 20044 56420 20100 56476
rect 50556 56420 50612 56476
rect 50660 56420 50716 56476
rect 50764 56420 50820 56476
rect 4476 55636 4532 55692
rect 4580 55636 4636 55692
rect 4684 55636 4740 55692
rect 35196 55636 35252 55692
rect 35300 55636 35356 55692
rect 35404 55636 35460 55692
rect 19836 54852 19892 54908
rect 19940 54852 19996 54908
rect 20044 54852 20100 54908
rect 50556 54852 50612 54908
rect 50660 54852 50716 54908
rect 50764 54852 50820 54908
rect 4476 54068 4532 54124
rect 4580 54068 4636 54124
rect 4684 54068 4740 54124
rect 35196 54068 35252 54124
rect 35300 54068 35356 54124
rect 35404 54068 35460 54124
rect 19836 53284 19892 53340
rect 19940 53284 19996 53340
rect 20044 53284 20100 53340
rect 50556 53284 50612 53340
rect 50660 53284 50716 53340
rect 50764 53284 50820 53340
rect 4476 52500 4532 52556
rect 4580 52500 4636 52556
rect 4684 52500 4740 52556
rect 35196 52500 35252 52556
rect 35300 52500 35356 52556
rect 35404 52500 35460 52556
rect 19836 51716 19892 51772
rect 19940 51716 19996 51772
rect 20044 51716 20100 51772
rect 50556 51716 50612 51772
rect 50660 51716 50716 51772
rect 50764 51716 50820 51772
rect 4476 50932 4532 50988
rect 4580 50932 4636 50988
rect 4684 50932 4740 50988
rect 35196 50932 35252 50988
rect 35300 50932 35356 50988
rect 35404 50932 35460 50988
rect 19836 50148 19892 50204
rect 19940 50148 19996 50204
rect 20044 50148 20100 50204
rect 50556 50148 50612 50204
rect 50660 50148 50716 50204
rect 50764 50148 50820 50204
rect 4476 49364 4532 49420
rect 4580 49364 4636 49420
rect 4684 49364 4740 49420
rect 35196 49364 35252 49420
rect 35300 49364 35356 49420
rect 35404 49364 35460 49420
rect 19836 48580 19892 48636
rect 19940 48580 19996 48636
rect 20044 48580 20100 48636
rect 19628 48300 19684 48356
rect 4476 47796 4532 47852
rect 4580 47796 4636 47852
rect 4684 47796 4740 47852
rect 50556 48580 50612 48636
rect 50660 48580 50716 48636
rect 50764 48580 50820 48636
rect 35196 47796 35252 47852
rect 35300 47796 35356 47852
rect 35404 47796 35460 47852
rect 19836 47012 19892 47068
rect 19940 47012 19996 47068
rect 20044 47012 20100 47068
rect 50556 47012 50612 47068
rect 50660 47012 50716 47068
rect 50764 47012 50820 47068
rect 12908 46844 12964 46900
rect 4476 46228 4532 46284
rect 4580 46228 4636 46284
rect 4684 46228 4740 46284
rect 35196 46228 35252 46284
rect 35300 46228 35356 46284
rect 35404 46228 35460 46284
rect 23660 46060 23716 46116
rect 26796 45836 26852 45892
rect 10556 45612 10612 45668
rect 18844 45500 18900 45556
rect 19836 45444 19892 45500
rect 19940 45444 19996 45500
rect 20044 45444 20100 45500
rect 50556 45444 50612 45500
rect 50660 45444 50716 45500
rect 50764 45444 50820 45500
rect 19292 44828 19348 44884
rect 4476 44660 4532 44716
rect 4580 44660 4636 44716
rect 4684 44660 4740 44716
rect 35196 44660 35252 44716
rect 35300 44660 35356 44716
rect 35404 44660 35460 44716
rect 18844 44604 18900 44660
rect 23212 44604 23268 44660
rect 26236 44380 26292 44436
rect 18060 44268 18116 44324
rect 16940 44156 16996 44212
rect 19836 43876 19892 43932
rect 19940 43876 19996 43932
rect 20044 43876 20100 43932
rect 50556 43876 50612 43932
rect 50660 43876 50716 43932
rect 50764 43876 50820 43932
rect 12124 43372 12180 43428
rect 23100 43372 23156 43428
rect 4476 43092 4532 43148
rect 4580 43092 4636 43148
rect 4684 43092 4740 43148
rect 35196 43092 35252 43148
rect 35300 43092 35356 43148
rect 35404 43092 35460 43148
rect 23884 42812 23940 42868
rect 10220 42476 10276 42532
rect 21868 42364 21924 42420
rect 23884 42364 23940 42420
rect 19836 42308 19892 42364
rect 19940 42308 19996 42364
rect 20044 42308 20100 42364
rect 50556 42308 50612 42364
rect 50660 42308 50716 42364
rect 50764 42308 50820 42364
rect 19292 41580 19348 41636
rect 4476 41524 4532 41580
rect 4580 41524 4636 41580
rect 4684 41524 4740 41580
rect 35196 41524 35252 41580
rect 35300 41524 35356 41580
rect 35404 41524 35460 41580
rect 21756 41132 21812 41188
rect 19836 40740 19892 40796
rect 19940 40740 19996 40796
rect 20044 40740 20100 40796
rect 50556 40740 50612 40796
rect 50660 40740 50716 40796
rect 50764 40740 50820 40796
rect 6636 40572 6692 40628
rect 18956 40460 19012 40516
rect 26124 40460 26180 40516
rect 11452 40348 11508 40404
rect 17724 40348 17780 40404
rect 21532 40124 21588 40180
rect 4476 39956 4532 40012
rect 4580 39956 4636 40012
rect 4684 39956 4740 40012
rect 35196 39956 35252 40012
rect 35300 39956 35356 40012
rect 35404 39956 35460 40012
rect 26124 39564 26180 39620
rect 23660 39452 23716 39508
rect 11788 39340 11844 39396
rect 19836 39172 19892 39228
rect 19940 39172 19996 39228
rect 20044 39172 20100 39228
rect 50556 39172 50612 39228
rect 50660 39172 50716 39228
rect 50764 39172 50820 39228
rect 16268 38892 16324 38948
rect 18172 38892 18228 38948
rect 15036 38668 15092 38724
rect 23212 38668 23268 38724
rect 4476 38388 4532 38444
rect 4580 38388 4636 38444
rect 4684 38388 4740 38444
rect 35196 38388 35252 38444
rect 35300 38388 35356 38444
rect 35404 38388 35460 38444
rect 16380 38220 16436 38276
rect 16604 38220 16660 38276
rect 21644 38220 21700 38276
rect 26236 38108 26292 38164
rect 15036 37996 15092 38052
rect 15484 37772 15540 37828
rect 19180 37660 19236 37716
rect 19836 37604 19892 37660
rect 19940 37604 19996 37660
rect 20044 37604 20100 37660
rect 50556 37604 50612 37660
rect 50660 37604 50716 37660
rect 50764 37604 50820 37660
rect 18284 37548 18340 37604
rect 26796 37436 26852 37492
rect 12908 37212 12964 37268
rect 18396 37212 18452 37268
rect 28028 37212 28084 37268
rect 19180 36876 19236 36932
rect 4476 36820 4532 36876
rect 4580 36820 4636 36876
rect 4684 36820 4740 36876
rect 15036 36764 15092 36820
rect 3164 36540 3220 36596
rect 11452 36540 11508 36596
rect 35196 36820 35252 36876
rect 35300 36820 35356 36876
rect 35404 36820 35460 36876
rect 14924 36204 14980 36260
rect 18396 36204 18452 36260
rect 21868 36204 21924 36260
rect 2828 36092 2884 36148
rect 15148 36092 15204 36148
rect 17724 36092 17780 36148
rect 18284 36092 18340 36148
rect 19292 36092 19348 36148
rect 28028 36092 28084 36148
rect 19836 36036 19892 36092
rect 19940 36036 19996 36092
rect 20044 36036 20100 36092
rect 50556 36036 50612 36092
rect 50660 36036 50716 36092
rect 50764 36036 50820 36092
rect 18844 35756 18900 35812
rect 20300 35644 20356 35700
rect 27804 35644 27860 35700
rect 2828 35532 2884 35588
rect 10220 35420 10276 35476
rect 10556 35420 10612 35476
rect 9884 35308 9940 35364
rect 10444 35308 10500 35364
rect 17052 35308 17108 35364
rect 18956 35308 19012 35364
rect 4476 35252 4532 35308
rect 4580 35252 4636 35308
rect 4684 35252 4740 35308
rect 35196 35252 35252 35308
rect 35300 35252 35356 35308
rect 35404 35252 35460 35308
rect 18844 35196 18900 35252
rect 18508 35084 18564 35140
rect 19404 35084 19460 35140
rect 10444 34972 10500 35028
rect 14476 34860 14532 34916
rect 16940 34860 16996 34916
rect 3164 34524 3220 34580
rect 19836 34468 19892 34524
rect 19940 34468 19996 34524
rect 20044 34468 20100 34524
rect 50556 34468 50612 34524
rect 50660 34468 50716 34524
rect 50764 34468 50820 34524
rect 14364 34412 14420 34468
rect 17612 34300 17668 34356
rect 21644 34300 21700 34356
rect 20300 33964 20356 34020
rect 21868 33964 21924 34020
rect 4476 33684 4532 33740
rect 4580 33684 4636 33740
rect 4684 33684 4740 33740
rect 6636 33516 6692 33572
rect 35196 33684 35252 33740
rect 35300 33684 35356 33740
rect 35404 33684 35460 33740
rect 13244 33404 13300 33460
rect 16380 33180 16436 33236
rect 19404 33068 19460 33124
rect 18172 32956 18228 33012
rect 19836 32900 19892 32956
rect 19940 32900 19996 32956
rect 20044 32900 20100 32956
rect 50556 32900 50612 32956
rect 50660 32900 50716 32956
rect 50764 32900 50820 32956
rect 20188 32844 20244 32900
rect 11900 32732 11956 32788
rect 10444 32508 10500 32564
rect 4476 32116 4532 32172
rect 4580 32116 4636 32172
rect 4684 32116 4740 32172
rect 35196 32116 35252 32172
rect 35300 32116 35356 32172
rect 35404 32116 35460 32172
rect 17612 31948 17668 32004
rect 20300 31836 20356 31892
rect 17052 31500 17108 31556
rect 18844 31388 18900 31444
rect 19836 31332 19892 31388
rect 19940 31332 19996 31388
rect 20044 31332 20100 31388
rect 50556 31332 50612 31388
rect 50660 31332 50716 31388
rect 50764 31332 50820 31388
rect 25900 31276 25956 31332
rect 5964 31164 6020 31220
rect 15036 31164 15092 31220
rect 18060 31164 18116 31220
rect 18732 31164 18788 31220
rect 14252 31052 14308 31108
rect 14476 31052 14532 31108
rect 11116 30940 11172 30996
rect 14924 30716 14980 30772
rect 4476 30548 4532 30604
rect 4580 30548 4636 30604
rect 4684 30548 4740 30604
rect 35196 30548 35252 30604
rect 35300 30548 35356 30604
rect 35404 30548 35460 30604
rect 11452 30492 11508 30548
rect 16268 30492 16324 30548
rect 21756 30380 21812 30436
rect 25900 30380 25956 30436
rect 14364 30268 14420 30324
rect 18732 30156 18788 30212
rect 28028 30156 28084 30212
rect 14924 30044 14980 30100
rect 20300 30044 20356 30100
rect 5740 29932 5796 29988
rect 11116 29932 11172 29988
rect 15148 29932 15204 29988
rect 11900 29708 11956 29764
rect 19836 29764 19892 29820
rect 19940 29764 19996 29820
rect 20044 29764 20100 29820
rect 5740 29372 5796 29428
rect 18732 29372 18788 29428
rect 50556 29764 50612 29820
rect 50660 29764 50716 29820
rect 50764 29764 50820 29820
rect 12684 29260 12740 29316
rect 14252 29148 14308 29204
rect 4476 28980 4532 29036
rect 4580 28980 4636 29036
rect 4684 28980 4740 29036
rect 35196 28980 35252 29036
rect 35300 28980 35356 29036
rect 35404 28980 35460 29036
rect 19404 28812 19460 28868
rect 14364 28700 14420 28756
rect 8652 28588 8708 28644
rect 19628 28364 19684 28420
rect 19836 28196 19892 28252
rect 19940 28196 19996 28252
rect 20044 28196 20100 28252
rect 50556 28196 50612 28252
rect 50660 28196 50716 28252
rect 50764 28196 50820 28252
rect 15036 28028 15092 28084
rect 12124 27804 12180 27860
rect 15036 27804 15092 27860
rect 8652 27692 8708 27748
rect 14252 27468 14308 27524
rect 4476 27412 4532 27468
rect 4580 27412 4636 27468
rect 4684 27412 4740 27468
rect 35196 27412 35252 27468
rect 35300 27412 35356 27468
rect 35404 27412 35460 27468
rect 21980 27132 22036 27188
rect 5964 27020 6020 27076
rect 11676 27020 11732 27076
rect 5740 26908 5796 26964
rect 11788 26796 11844 26852
rect 12684 26684 12740 26740
rect 11452 26572 11508 26628
rect 13244 26460 13300 26516
rect 19836 26628 19892 26684
rect 19940 26628 19996 26684
rect 20044 26628 20100 26684
rect 50556 26628 50612 26684
rect 50660 26628 50716 26684
rect 50764 26628 50820 26684
rect 20188 26572 20244 26628
rect 4476 25844 4532 25900
rect 4580 25844 4636 25900
rect 4684 25844 4740 25900
rect 35196 25844 35252 25900
rect 35300 25844 35356 25900
rect 35404 25844 35460 25900
rect 14924 25788 14980 25844
rect 19404 25452 19460 25508
rect 20188 25340 20244 25396
rect 11676 25228 11732 25284
rect 19836 25060 19892 25116
rect 19940 25060 19996 25116
rect 20044 25060 20100 25116
rect 50556 25060 50612 25116
rect 50660 25060 50716 25116
rect 50764 25060 50820 25116
rect 18508 24556 18564 24612
rect 4476 24276 4532 24332
rect 4580 24276 4636 24332
rect 4684 24276 4740 24332
rect 35196 24276 35252 24332
rect 35300 24276 35356 24332
rect 35404 24276 35460 24332
rect 15484 23884 15540 23940
rect 21532 23772 21588 23828
rect 19836 23492 19892 23548
rect 19940 23492 19996 23548
rect 20044 23492 20100 23548
rect 50556 23492 50612 23548
rect 50660 23492 50716 23548
rect 50764 23492 50820 23548
rect 4476 22708 4532 22764
rect 4580 22708 4636 22764
rect 4684 22708 4740 22764
rect 35196 22708 35252 22764
rect 35300 22708 35356 22764
rect 35404 22708 35460 22764
rect 19836 21924 19892 21980
rect 19940 21924 19996 21980
rect 20044 21924 20100 21980
rect 50556 21924 50612 21980
rect 50660 21924 50716 21980
rect 50764 21924 50820 21980
rect 23100 21756 23156 21812
rect 27804 21644 27860 21700
rect 4476 21140 4532 21196
rect 4580 21140 4636 21196
rect 4684 21140 4740 21196
rect 35196 21140 35252 21196
rect 35300 21140 35356 21196
rect 35404 21140 35460 21196
rect 19836 20356 19892 20412
rect 19940 20356 19996 20412
rect 20044 20356 20100 20412
rect 50556 20356 50612 20412
rect 50660 20356 50716 20412
rect 50764 20356 50820 20412
rect 4476 19572 4532 19628
rect 4580 19572 4636 19628
rect 4684 19572 4740 19628
rect 35196 19572 35252 19628
rect 35300 19572 35356 19628
rect 35404 19572 35460 19628
rect 19836 18788 19892 18844
rect 19940 18788 19996 18844
rect 20044 18788 20100 18844
rect 50556 18788 50612 18844
rect 50660 18788 50716 18844
rect 50764 18788 50820 18844
rect 4476 18004 4532 18060
rect 4580 18004 4636 18060
rect 4684 18004 4740 18060
rect 35196 18004 35252 18060
rect 35300 18004 35356 18060
rect 35404 18004 35460 18060
rect 19836 17220 19892 17276
rect 19940 17220 19996 17276
rect 20044 17220 20100 17276
rect 50556 17220 50612 17276
rect 50660 17220 50716 17276
rect 50764 17220 50820 17276
rect 4476 16436 4532 16492
rect 4580 16436 4636 16492
rect 4684 16436 4740 16492
rect 35196 16436 35252 16492
rect 35300 16436 35356 16492
rect 35404 16436 35460 16492
rect 19836 15652 19892 15708
rect 19940 15652 19996 15708
rect 20044 15652 20100 15708
rect 50556 15652 50612 15708
rect 50660 15652 50716 15708
rect 50764 15652 50820 15708
rect 4476 14868 4532 14924
rect 4580 14868 4636 14924
rect 4684 14868 4740 14924
rect 35196 14868 35252 14924
rect 35300 14868 35356 14924
rect 35404 14868 35460 14924
rect 19836 14084 19892 14140
rect 19940 14084 19996 14140
rect 20044 14084 20100 14140
rect 50556 14084 50612 14140
rect 50660 14084 50716 14140
rect 50764 14084 50820 14140
rect 4476 13300 4532 13356
rect 4580 13300 4636 13356
rect 4684 13300 4740 13356
rect 35196 13300 35252 13356
rect 35300 13300 35356 13356
rect 35404 13300 35460 13356
rect 19836 12516 19892 12572
rect 19940 12516 19996 12572
rect 20044 12516 20100 12572
rect 50556 12516 50612 12572
rect 50660 12516 50716 12572
rect 50764 12516 50820 12572
rect 4476 11732 4532 11788
rect 4580 11732 4636 11788
rect 4684 11732 4740 11788
rect 35196 11732 35252 11788
rect 35300 11732 35356 11788
rect 35404 11732 35460 11788
rect 19836 10948 19892 11004
rect 19940 10948 19996 11004
rect 20044 10948 20100 11004
rect 50556 10948 50612 11004
rect 50660 10948 50716 11004
rect 50764 10948 50820 11004
rect 4476 10164 4532 10220
rect 4580 10164 4636 10220
rect 4684 10164 4740 10220
rect 35196 10164 35252 10220
rect 35300 10164 35356 10220
rect 35404 10164 35460 10220
rect 19836 9380 19892 9436
rect 19940 9380 19996 9436
rect 20044 9380 20100 9436
rect 50556 9380 50612 9436
rect 50660 9380 50716 9436
rect 50764 9380 50820 9436
rect 4476 8596 4532 8652
rect 4580 8596 4636 8652
rect 4684 8596 4740 8652
rect 35196 8596 35252 8652
rect 35300 8596 35356 8652
rect 35404 8596 35460 8652
rect 19836 7812 19892 7868
rect 19940 7812 19996 7868
rect 20044 7812 20100 7868
rect 50556 7812 50612 7868
rect 50660 7812 50716 7868
rect 50764 7812 50820 7868
rect 4476 7028 4532 7084
rect 4580 7028 4636 7084
rect 4684 7028 4740 7084
rect 35196 7028 35252 7084
rect 35300 7028 35356 7084
rect 35404 7028 35460 7084
rect 19836 6244 19892 6300
rect 19940 6244 19996 6300
rect 20044 6244 20100 6300
rect 50556 6244 50612 6300
rect 50660 6244 50716 6300
rect 50764 6244 50820 6300
rect 4476 5460 4532 5516
rect 4580 5460 4636 5516
rect 4684 5460 4740 5516
rect 35196 5460 35252 5516
rect 35300 5460 35356 5516
rect 35404 5460 35460 5516
rect 19836 4676 19892 4732
rect 19940 4676 19996 4732
rect 20044 4676 20100 4732
rect 50556 4676 50612 4732
rect 50660 4676 50716 4732
rect 50764 4676 50820 4732
rect 4476 3892 4532 3948
rect 4580 3892 4636 3948
rect 4684 3892 4740 3948
rect 35196 3892 35252 3948
rect 35300 3892 35356 3948
rect 35404 3892 35460 3948
rect 19836 3108 19892 3164
rect 19940 3108 19996 3164
rect 20044 3108 20100 3164
rect 50556 3108 50612 3164
rect 50660 3108 50716 3164
rect 50764 3108 50820 3164
<< metal4 >>
rect 4448 55692 4768 56508
rect 4448 55636 4476 55692
rect 4532 55636 4580 55692
rect 4636 55636 4684 55692
rect 4740 55636 4768 55692
rect 4448 54124 4768 55636
rect 4448 54068 4476 54124
rect 4532 54068 4580 54124
rect 4636 54068 4684 54124
rect 4740 54068 4768 54124
rect 4448 52556 4768 54068
rect 4448 52500 4476 52556
rect 4532 52500 4580 52556
rect 4636 52500 4684 52556
rect 4740 52500 4768 52556
rect 4448 50988 4768 52500
rect 4448 50932 4476 50988
rect 4532 50932 4580 50988
rect 4636 50932 4684 50988
rect 4740 50932 4768 50988
rect 4448 49420 4768 50932
rect 4448 49364 4476 49420
rect 4532 49364 4580 49420
rect 4636 49364 4684 49420
rect 4740 49364 4768 49420
rect 4448 47852 4768 49364
rect 19808 56476 20128 56508
rect 19808 56420 19836 56476
rect 19892 56420 19940 56476
rect 19996 56420 20044 56476
rect 20100 56420 20128 56476
rect 19808 54908 20128 56420
rect 19808 54852 19836 54908
rect 19892 54852 19940 54908
rect 19996 54852 20044 54908
rect 20100 54852 20128 54908
rect 19808 53340 20128 54852
rect 19808 53284 19836 53340
rect 19892 53284 19940 53340
rect 19996 53284 20044 53340
rect 20100 53284 20128 53340
rect 19808 51772 20128 53284
rect 19808 51716 19836 51772
rect 19892 51716 19940 51772
rect 19996 51716 20044 51772
rect 20100 51716 20128 51772
rect 19808 50204 20128 51716
rect 19808 50148 19836 50204
rect 19892 50148 19940 50204
rect 19996 50148 20044 50204
rect 20100 50148 20128 50204
rect 19808 48636 20128 50148
rect 19808 48580 19836 48636
rect 19892 48580 19940 48636
rect 19996 48580 20044 48636
rect 20100 48580 20128 48636
rect 4448 47796 4476 47852
rect 4532 47796 4580 47852
rect 4636 47796 4684 47852
rect 4740 47796 4768 47852
rect 4448 46284 4768 47796
rect 19628 48356 19684 48366
rect 4448 46228 4476 46284
rect 4532 46228 4580 46284
rect 4636 46228 4684 46284
rect 4740 46228 4768 46284
rect 4448 44716 4768 46228
rect 12908 46900 12964 46910
rect 4448 44660 4476 44716
rect 4532 44660 4580 44716
rect 4636 44660 4684 44716
rect 4740 44660 4768 44716
rect 4448 43148 4768 44660
rect 4448 43092 4476 43148
rect 4532 43092 4580 43148
rect 4636 43092 4684 43148
rect 4740 43092 4768 43148
rect 4448 41580 4768 43092
rect 10556 45668 10612 45678
rect 4448 41524 4476 41580
rect 4532 41524 4580 41580
rect 4636 41524 4684 41580
rect 4740 41524 4768 41580
rect 4448 40012 4768 41524
rect 10220 42532 10276 42542
rect 4448 39956 4476 40012
rect 4532 39956 4580 40012
rect 4636 39956 4684 40012
rect 4740 39956 4768 40012
rect 4448 38444 4768 39956
rect 4448 38388 4476 38444
rect 4532 38388 4580 38444
rect 4636 38388 4684 38444
rect 4740 38388 4768 38444
rect 4448 36876 4768 38388
rect 4448 36820 4476 36876
rect 4532 36820 4580 36876
rect 4636 36820 4684 36876
rect 4740 36820 4768 36876
rect 3164 36596 3220 36606
rect 2828 36148 2884 36158
rect 2828 35588 2884 36092
rect 2828 35522 2884 35532
rect 3164 34580 3220 36540
rect 3164 34514 3220 34524
rect 4448 35308 4768 36820
rect 4448 35252 4476 35308
rect 4532 35252 4580 35308
rect 4636 35252 4684 35308
rect 4740 35252 4768 35308
rect 4448 33740 4768 35252
rect 4448 33684 4476 33740
rect 4532 33684 4580 33740
rect 4636 33684 4684 33740
rect 4740 33684 4768 33740
rect 4448 32172 4768 33684
rect 6636 40628 6692 40638
rect 6636 33572 6692 40572
rect 10220 35476 10276 42476
rect 10220 35410 10276 35420
rect 10556 35476 10612 45612
rect 12124 43428 12180 43438
rect 11452 40404 11508 40414
rect 11452 36596 11508 40348
rect 11452 36530 11508 36540
rect 11788 39396 11844 39406
rect 10556 35410 10612 35420
rect 9884 35364 9940 35374
rect 10444 35364 10500 35374
rect 9884 35252 10500 35308
rect 6636 33506 6692 33516
rect 10444 35028 10500 35038
rect 10444 32564 10500 34972
rect 10444 32498 10500 32508
rect 4448 32116 4476 32172
rect 4532 32116 4580 32172
rect 4636 32116 4684 32172
rect 4740 32116 4768 32172
rect 4448 30604 4768 32116
rect 4448 30548 4476 30604
rect 4532 30548 4580 30604
rect 4636 30548 4684 30604
rect 4740 30548 4768 30604
rect 4448 29036 4768 30548
rect 5964 31220 6020 31230
rect 4448 28980 4476 29036
rect 4532 28980 4580 29036
rect 4636 28980 4684 29036
rect 4740 28980 4768 29036
rect 4448 27468 4768 28980
rect 4448 27412 4476 27468
rect 4532 27412 4580 27468
rect 4636 27412 4684 27468
rect 4740 27412 4768 27468
rect 4448 25900 4768 27412
rect 5740 29988 5796 29998
rect 5740 29428 5796 29932
rect 5740 26964 5796 29372
rect 5964 27076 6020 31164
rect 11116 30996 11172 31006
rect 11116 29988 11172 30940
rect 11116 29922 11172 29932
rect 11452 30548 11508 30558
rect 8652 28644 8708 28654
rect 8652 27748 8708 28588
rect 8652 27682 8708 27692
rect 5964 27010 6020 27020
rect 5740 26898 5796 26908
rect 11452 26628 11508 30492
rect 11452 26562 11508 26572
rect 11676 27076 11732 27086
rect 4448 25844 4476 25900
rect 4532 25844 4580 25900
rect 4636 25844 4684 25900
rect 4740 25844 4768 25900
rect 4448 24332 4768 25844
rect 11676 25284 11732 27020
rect 11788 26852 11844 39340
rect 11900 32788 11956 32798
rect 11900 29764 11956 32732
rect 11900 29698 11956 29708
rect 12124 27860 12180 43372
rect 12908 37268 12964 46844
rect 18844 45556 18900 45566
rect 18844 44660 18900 45500
rect 18060 44324 18116 44334
rect 16940 44212 16996 44222
rect 16268 38948 16324 38958
rect 15036 38724 15092 38734
rect 15036 38052 15092 38668
rect 15036 37986 15092 37996
rect 16268 38458 16324 38892
rect 16268 38402 16660 38458
rect 12908 37202 12964 37212
rect 15484 37828 15540 37838
rect 15036 36820 15092 36830
rect 14924 36260 14980 36270
rect 14476 34916 14532 34926
rect 14364 34468 14420 34478
rect 13244 33460 13300 33470
rect 12124 27794 12180 27804
rect 12684 29316 12740 29326
rect 11788 26786 11844 26796
rect 12684 26740 12740 29260
rect 12684 26674 12740 26684
rect 13244 26516 13300 33404
rect 14252 31108 14308 31118
rect 14252 29204 14308 31052
rect 14252 27524 14308 29148
rect 14364 30324 14420 34412
rect 14476 31108 14532 34860
rect 14476 31042 14532 31052
rect 14924 30772 14980 36204
rect 14924 30706 14980 30716
rect 15036 31220 15092 36764
rect 14364 28756 14420 30268
rect 14364 28690 14420 28700
rect 14924 30100 14980 30110
rect 14252 27458 14308 27468
rect 13244 26450 13300 26460
rect 14924 25844 14980 30044
rect 15036 28084 15092 31164
rect 15148 36148 15204 36158
rect 15148 29988 15204 36092
rect 15148 29922 15204 29932
rect 15036 27860 15092 28028
rect 15036 27794 15092 27804
rect 14924 25778 14980 25788
rect 11676 25218 11732 25228
rect 4448 24276 4476 24332
rect 4532 24276 4580 24332
rect 4636 24276 4684 24332
rect 4740 24276 4768 24332
rect 4448 22764 4768 24276
rect 15484 23940 15540 37772
rect 16268 30548 16324 38402
rect 16380 38276 16436 38286
rect 16380 33236 16436 38220
rect 16604 38276 16660 38402
rect 16604 38210 16660 38220
rect 16940 34916 16996 44156
rect 17724 40404 17780 40414
rect 17724 36148 17780 40348
rect 17724 36082 17780 36092
rect 16940 34850 16996 34860
rect 17052 35364 17108 35374
rect 16380 33170 16436 33180
rect 17052 31556 17108 35308
rect 17612 34356 17668 34366
rect 17612 32004 17668 34300
rect 17612 31938 17668 31948
rect 17052 31490 17108 31500
rect 18060 31220 18116 44268
rect 18172 38948 18228 38958
rect 18172 33012 18228 38892
rect 18284 37604 18340 37614
rect 18284 36148 18340 37548
rect 18396 37268 18452 37278
rect 18396 36260 18452 37212
rect 18396 36194 18452 36204
rect 18284 36082 18340 36092
rect 18844 35812 18900 44604
rect 19292 44884 19348 44894
rect 19292 41636 19348 44828
rect 18844 35746 18900 35756
rect 18956 40516 19012 40526
rect 18956 35364 19012 40460
rect 19180 37716 19236 37726
rect 19180 36932 19236 37660
rect 19180 36866 19236 36876
rect 19292 36148 19348 41580
rect 19292 36082 19348 36092
rect 18956 35298 19012 35308
rect 18844 35252 18900 35262
rect 18172 32946 18228 32956
rect 18508 35140 18564 35150
rect 18060 31154 18116 31164
rect 16268 30482 16324 30492
rect 18508 24612 18564 35084
rect 18844 31444 18900 35196
rect 18844 31378 18900 31388
rect 19404 35140 19460 35150
rect 19404 33124 19460 35084
rect 18732 31220 18788 31230
rect 18732 30212 18788 31164
rect 18732 29428 18788 30156
rect 18732 29362 18788 29372
rect 19404 28868 19460 33068
rect 19404 25508 19460 28812
rect 19628 28420 19684 48300
rect 19628 28354 19684 28364
rect 19808 47068 20128 48580
rect 19808 47012 19836 47068
rect 19892 47012 19940 47068
rect 19996 47012 20044 47068
rect 20100 47012 20128 47068
rect 19808 45500 20128 47012
rect 35168 55692 35488 56508
rect 35168 55636 35196 55692
rect 35252 55636 35300 55692
rect 35356 55636 35404 55692
rect 35460 55636 35488 55692
rect 35168 54124 35488 55636
rect 35168 54068 35196 54124
rect 35252 54068 35300 54124
rect 35356 54068 35404 54124
rect 35460 54068 35488 54124
rect 35168 52556 35488 54068
rect 35168 52500 35196 52556
rect 35252 52500 35300 52556
rect 35356 52500 35404 52556
rect 35460 52500 35488 52556
rect 35168 50988 35488 52500
rect 35168 50932 35196 50988
rect 35252 50932 35300 50988
rect 35356 50932 35404 50988
rect 35460 50932 35488 50988
rect 35168 49420 35488 50932
rect 35168 49364 35196 49420
rect 35252 49364 35300 49420
rect 35356 49364 35404 49420
rect 35460 49364 35488 49420
rect 35168 47852 35488 49364
rect 35168 47796 35196 47852
rect 35252 47796 35300 47852
rect 35356 47796 35404 47852
rect 35460 47796 35488 47852
rect 35168 46284 35488 47796
rect 35168 46228 35196 46284
rect 35252 46228 35300 46284
rect 35356 46228 35404 46284
rect 35460 46228 35488 46284
rect 19808 45444 19836 45500
rect 19892 45444 19940 45500
rect 19996 45444 20044 45500
rect 20100 45444 20128 45500
rect 19808 43932 20128 45444
rect 23660 46116 23716 46126
rect 19808 43876 19836 43932
rect 19892 43876 19940 43932
rect 19996 43876 20044 43932
rect 20100 43876 20128 43932
rect 19808 42364 20128 43876
rect 23212 44660 23268 44670
rect 23100 43428 23156 43438
rect 19808 42308 19836 42364
rect 19892 42308 19940 42364
rect 19996 42308 20044 42364
rect 20100 42308 20128 42364
rect 19808 40796 20128 42308
rect 21868 42420 21924 42430
rect 19808 40740 19836 40796
rect 19892 40740 19940 40796
rect 19996 40740 20044 40796
rect 20100 40740 20128 40796
rect 19808 39228 20128 40740
rect 21756 41188 21812 41198
rect 19808 39172 19836 39228
rect 19892 39172 19940 39228
rect 19996 39172 20044 39228
rect 20100 39172 20128 39228
rect 19808 37660 20128 39172
rect 19808 37604 19836 37660
rect 19892 37604 19940 37660
rect 19996 37604 20044 37660
rect 20100 37604 20128 37660
rect 19808 36092 20128 37604
rect 19808 36036 19836 36092
rect 19892 36036 19940 36092
rect 19996 36036 20044 36092
rect 20100 36036 20128 36092
rect 19808 34524 20128 36036
rect 21532 40180 21588 40190
rect 19808 34468 19836 34524
rect 19892 34468 19940 34524
rect 19996 34468 20044 34524
rect 20100 34468 20128 34524
rect 19808 32956 20128 34468
rect 20300 35700 20356 35710
rect 20300 34020 20356 35644
rect 20300 33954 20356 33964
rect 19808 32900 19836 32956
rect 19892 32900 19940 32956
rect 19996 32900 20044 32956
rect 20100 32900 20128 32956
rect 19808 31388 20128 32900
rect 19808 31332 19836 31388
rect 19892 31332 19940 31388
rect 19996 31332 20044 31388
rect 20100 31332 20128 31388
rect 19808 29820 20128 31332
rect 19808 29764 19836 29820
rect 19892 29764 19940 29820
rect 19996 29764 20044 29820
rect 20100 29764 20128 29820
rect 19404 25442 19460 25452
rect 19808 28252 20128 29764
rect 19808 28196 19836 28252
rect 19892 28196 19940 28252
rect 19996 28196 20044 28252
rect 20100 28196 20128 28252
rect 19808 26684 20128 28196
rect 19808 26628 19836 26684
rect 19892 26628 19940 26684
rect 19996 26628 20044 26684
rect 20100 26628 20128 26684
rect 18508 24546 18564 24556
rect 19808 25116 20128 26628
rect 20188 32900 20244 32910
rect 20188 26628 20244 32844
rect 20300 31892 20356 31902
rect 20300 30100 20356 31836
rect 20300 30034 20356 30044
rect 20188 25396 20244 26572
rect 20188 25330 20244 25340
rect 19808 25060 19836 25116
rect 19892 25060 19940 25116
rect 19996 25060 20044 25116
rect 20100 25060 20128 25116
rect 15484 23874 15540 23884
rect 4448 22708 4476 22764
rect 4532 22708 4580 22764
rect 4636 22708 4684 22764
rect 4740 22708 4768 22764
rect 4448 21196 4768 22708
rect 4448 21140 4476 21196
rect 4532 21140 4580 21196
rect 4636 21140 4684 21196
rect 4740 21140 4768 21196
rect 4448 19628 4768 21140
rect 4448 19572 4476 19628
rect 4532 19572 4580 19628
rect 4636 19572 4684 19628
rect 4740 19572 4768 19628
rect 4448 18060 4768 19572
rect 4448 18004 4476 18060
rect 4532 18004 4580 18060
rect 4636 18004 4684 18060
rect 4740 18004 4768 18060
rect 4448 16492 4768 18004
rect 4448 16436 4476 16492
rect 4532 16436 4580 16492
rect 4636 16436 4684 16492
rect 4740 16436 4768 16492
rect 4448 14924 4768 16436
rect 4448 14868 4476 14924
rect 4532 14868 4580 14924
rect 4636 14868 4684 14924
rect 4740 14868 4768 14924
rect 4448 13356 4768 14868
rect 4448 13300 4476 13356
rect 4532 13300 4580 13356
rect 4636 13300 4684 13356
rect 4740 13300 4768 13356
rect 4448 11788 4768 13300
rect 4448 11732 4476 11788
rect 4532 11732 4580 11788
rect 4636 11732 4684 11788
rect 4740 11732 4768 11788
rect 4448 10220 4768 11732
rect 4448 10164 4476 10220
rect 4532 10164 4580 10220
rect 4636 10164 4684 10220
rect 4740 10164 4768 10220
rect 4448 8652 4768 10164
rect 4448 8596 4476 8652
rect 4532 8596 4580 8652
rect 4636 8596 4684 8652
rect 4740 8596 4768 8652
rect 4448 7084 4768 8596
rect 4448 7028 4476 7084
rect 4532 7028 4580 7084
rect 4636 7028 4684 7084
rect 4740 7028 4768 7084
rect 4448 5516 4768 7028
rect 4448 5460 4476 5516
rect 4532 5460 4580 5516
rect 4636 5460 4684 5516
rect 4740 5460 4768 5516
rect 4448 3948 4768 5460
rect 4448 3892 4476 3948
rect 4532 3892 4580 3948
rect 4636 3892 4684 3948
rect 4740 3892 4768 3948
rect 4448 3076 4768 3892
rect 19808 23548 20128 25060
rect 21532 23828 21588 40124
rect 21644 38276 21700 38286
rect 21644 34356 21700 38220
rect 21644 34290 21700 34300
rect 21756 30436 21812 41132
rect 21868 38668 21924 42364
rect 21868 38612 22036 38668
rect 21868 36260 21924 36270
rect 21868 34020 21924 36204
rect 21868 33954 21924 33964
rect 21756 30370 21812 30380
rect 21980 27188 22036 38612
rect 21980 27122 22036 27132
rect 21532 23762 21588 23772
rect 19808 23492 19836 23548
rect 19892 23492 19940 23548
rect 19996 23492 20044 23548
rect 20100 23492 20128 23548
rect 19808 21980 20128 23492
rect 19808 21924 19836 21980
rect 19892 21924 19940 21980
rect 19996 21924 20044 21980
rect 20100 21924 20128 21980
rect 19808 20412 20128 21924
rect 23100 21812 23156 43372
rect 23212 38724 23268 44604
rect 23660 39508 23716 46060
rect 26796 45892 26852 45902
rect 26236 44436 26292 44446
rect 23884 42868 23940 42878
rect 23884 42420 23940 42812
rect 23884 42354 23940 42364
rect 26124 40516 26180 40526
rect 26124 39620 26180 40460
rect 26124 39554 26180 39564
rect 23660 39442 23716 39452
rect 23212 38658 23268 38668
rect 26236 38164 26292 44380
rect 26236 38098 26292 38108
rect 26796 37492 26852 45836
rect 26796 37426 26852 37436
rect 35168 44716 35488 46228
rect 35168 44660 35196 44716
rect 35252 44660 35300 44716
rect 35356 44660 35404 44716
rect 35460 44660 35488 44716
rect 35168 43148 35488 44660
rect 35168 43092 35196 43148
rect 35252 43092 35300 43148
rect 35356 43092 35404 43148
rect 35460 43092 35488 43148
rect 35168 41580 35488 43092
rect 35168 41524 35196 41580
rect 35252 41524 35300 41580
rect 35356 41524 35404 41580
rect 35460 41524 35488 41580
rect 35168 40012 35488 41524
rect 35168 39956 35196 40012
rect 35252 39956 35300 40012
rect 35356 39956 35404 40012
rect 35460 39956 35488 40012
rect 35168 38444 35488 39956
rect 35168 38388 35196 38444
rect 35252 38388 35300 38444
rect 35356 38388 35404 38444
rect 35460 38388 35488 38444
rect 28028 37268 28084 37278
rect 28028 36148 28084 37212
rect 27804 35700 27860 35710
rect 25900 31332 25956 31342
rect 25900 30436 25956 31276
rect 25900 30370 25956 30380
rect 23100 21746 23156 21756
rect 27804 21700 27860 35644
rect 28028 30212 28084 36092
rect 28028 30146 28084 30156
rect 35168 36876 35488 38388
rect 35168 36820 35196 36876
rect 35252 36820 35300 36876
rect 35356 36820 35404 36876
rect 35460 36820 35488 36876
rect 35168 35308 35488 36820
rect 35168 35252 35196 35308
rect 35252 35252 35300 35308
rect 35356 35252 35404 35308
rect 35460 35252 35488 35308
rect 35168 33740 35488 35252
rect 35168 33684 35196 33740
rect 35252 33684 35300 33740
rect 35356 33684 35404 33740
rect 35460 33684 35488 33740
rect 35168 32172 35488 33684
rect 35168 32116 35196 32172
rect 35252 32116 35300 32172
rect 35356 32116 35404 32172
rect 35460 32116 35488 32172
rect 35168 30604 35488 32116
rect 35168 30548 35196 30604
rect 35252 30548 35300 30604
rect 35356 30548 35404 30604
rect 35460 30548 35488 30604
rect 27804 21634 27860 21644
rect 35168 29036 35488 30548
rect 35168 28980 35196 29036
rect 35252 28980 35300 29036
rect 35356 28980 35404 29036
rect 35460 28980 35488 29036
rect 35168 27468 35488 28980
rect 35168 27412 35196 27468
rect 35252 27412 35300 27468
rect 35356 27412 35404 27468
rect 35460 27412 35488 27468
rect 35168 25900 35488 27412
rect 35168 25844 35196 25900
rect 35252 25844 35300 25900
rect 35356 25844 35404 25900
rect 35460 25844 35488 25900
rect 35168 24332 35488 25844
rect 35168 24276 35196 24332
rect 35252 24276 35300 24332
rect 35356 24276 35404 24332
rect 35460 24276 35488 24332
rect 35168 22764 35488 24276
rect 35168 22708 35196 22764
rect 35252 22708 35300 22764
rect 35356 22708 35404 22764
rect 35460 22708 35488 22764
rect 19808 20356 19836 20412
rect 19892 20356 19940 20412
rect 19996 20356 20044 20412
rect 20100 20356 20128 20412
rect 19808 18844 20128 20356
rect 19808 18788 19836 18844
rect 19892 18788 19940 18844
rect 19996 18788 20044 18844
rect 20100 18788 20128 18844
rect 19808 17276 20128 18788
rect 19808 17220 19836 17276
rect 19892 17220 19940 17276
rect 19996 17220 20044 17276
rect 20100 17220 20128 17276
rect 19808 15708 20128 17220
rect 19808 15652 19836 15708
rect 19892 15652 19940 15708
rect 19996 15652 20044 15708
rect 20100 15652 20128 15708
rect 19808 14140 20128 15652
rect 19808 14084 19836 14140
rect 19892 14084 19940 14140
rect 19996 14084 20044 14140
rect 20100 14084 20128 14140
rect 19808 12572 20128 14084
rect 19808 12516 19836 12572
rect 19892 12516 19940 12572
rect 19996 12516 20044 12572
rect 20100 12516 20128 12572
rect 19808 11004 20128 12516
rect 19808 10948 19836 11004
rect 19892 10948 19940 11004
rect 19996 10948 20044 11004
rect 20100 10948 20128 11004
rect 19808 9436 20128 10948
rect 19808 9380 19836 9436
rect 19892 9380 19940 9436
rect 19996 9380 20044 9436
rect 20100 9380 20128 9436
rect 19808 7868 20128 9380
rect 19808 7812 19836 7868
rect 19892 7812 19940 7868
rect 19996 7812 20044 7868
rect 20100 7812 20128 7868
rect 19808 6300 20128 7812
rect 19808 6244 19836 6300
rect 19892 6244 19940 6300
rect 19996 6244 20044 6300
rect 20100 6244 20128 6300
rect 19808 4732 20128 6244
rect 19808 4676 19836 4732
rect 19892 4676 19940 4732
rect 19996 4676 20044 4732
rect 20100 4676 20128 4732
rect 19808 3164 20128 4676
rect 19808 3108 19836 3164
rect 19892 3108 19940 3164
rect 19996 3108 20044 3164
rect 20100 3108 20128 3164
rect 19808 3076 20128 3108
rect 35168 21196 35488 22708
rect 35168 21140 35196 21196
rect 35252 21140 35300 21196
rect 35356 21140 35404 21196
rect 35460 21140 35488 21196
rect 35168 19628 35488 21140
rect 35168 19572 35196 19628
rect 35252 19572 35300 19628
rect 35356 19572 35404 19628
rect 35460 19572 35488 19628
rect 35168 18060 35488 19572
rect 35168 18004 35196 18060
rect 35252 18004 35300 18060
rect 35356 18004 35404 18060
rect 35460 18004 35488 18060
rect 35168 16492 35488 18004
rect 35168 16436 35196 16492
rect 35252 16436 35300 16492
rect 35356 16436 35404 16492
rect 35460 16436 35488 16492
rect 35168 14924 35488 16436
rect 35168 14868 35196 14924
rect 35252 14868 35300 14924
rect 35356 14868 35404 14924
rect 35460 14868 35488 14924
rect 35168 13356 35488 14868
rect 35168 13300 35196 13356
rect 35252 13300 35300 13356
rect 35356 13300 35404 13356
rect 35460 13300 35488 13356
rect 35168 11788 35488 13300
rect 35168 11732 35196 11788
rect 35252 11732 35300 11788
rect 35356 11732 35404 11788
rect 35460 11732 35488 11788
rect 35168 10220 35488 11732
rect 35168 10164 35196 10220
rect 35252 10164 35300 10220
rect 35356 10164 35404 10220
rect 35460 10164 35488 10220
rect 35168 8652 35488 10164
rect 35168 8596 35196 8652
rect 35252 8596 35300 8652
rect 35356 8596 35404 8652
rect 35460 8596 35488 8652
rect 35168 7084 35488 8596
rect 35168 7028 35196 7084
rect 35252 7028 35300 7084
rect 35356 7028 35404 7084
rect 35460 7028 35488 7084
rect 35168 5516 35488 7028
rect 35168 5460 35196 5516
rect 35252 5460 35300 5516
rect 35356 5460 35404 5516
rect 35460 5460 35488 5516
rect 35168 3948 35488 5460
rect 35168 3892 35196 3948
rect 35252 3892 35300 3948
rect 35356 3892 35404 3948
rect 35460 3892 35488 3948
rect 35168 3076 35488 3892
rect 50528 56476 50848 56508
rect 50528 56420 50556 56476
rect 50612 56420 50660 56476
rect 50716 56420 50764 56476
rect 50820 56420 50848 56476
rect 50528 54908 50848 56420
rect 50528 54852 50556 54908
rect 50612 54852 50660 54908
rect 50716 54852 50764 54908
rect 50820 54852 50848 54908
rect 50528 53340 50848 54852
rect 50528 53284 50556 53340
rect 50612 53284 50660 53340
rect 50716 53284 50764 53340
rect 50820 53284 50848 53340
rect 50528 51772 50848 53284
rect 50528 51716 50556 51772
rect 50612 51716 50660 51772
rect 50716 51716 50764 51772
rect 50820 51716 50848 51772
rect 50528 50204 50848 51716
rect 50528 50148 50556 50204
rect 50612 50148 50660 50204
rect 50716 50148 50764 50204
rect 50820 50148 50848 50204
rect 50528 48636 50848 50148
rect 50528 48580 50556 48636
rect 50612 48580 50660 48636
rect 50716 48580 50764 48636
rect 50820 48580 50848 48636
rect 50528 47068 50848 48580
rect 50528 47012 50556 47068
rect 50612 47012 50660 47068
rect 50716 47012 50764 47068
rect 50820 47012 50848 47068
rect 50528 45500 50848 47012
rect 50528 45444 50556 45500
rect 50612 45444 50660 45500
rect 50716 45444 50764 45500
rect 50820 45444 50848 45500
rect 50528 43932 50848 45444
rect 50528 43876 50556 43932
rect 50612 43876 50660 43932
rect 50716 43876 50764 43932
rect 50820 43876 50848 43932
rect 50528 42364 50848 43876
rect 50528 42308 50556 42364
rect 50612 42308 50660 42364
rect 50716 42308 50764 42364
rect 50820 42308 50848 42364
rect 50528 40796 50848 42308
rect 50528 40740 50556 40796
rect 50612 40740 50660 40796
rect 50716 40740 50764 40796
rect 50820 40740 50848 40796
rect 50528 39228 50848 40740
rect 50528 39172 50556 39228
rect 50612 39172 50660 39228
rect 50716 39172 50764 39228
rect 50820 39172 50848 39228
rect 50528 37660 50848 39172
rect 50528 37604 50556 37660
rect 50612 37604 50660 37660
rect 50716 37604 50764 37660
rect 50820 37604 50848 37660
rect 50528 36092 50848 37604
rect 50528 36036 50556 36092
rect 50612 36036 50660 36092
rect 50716 36036 50764 36092
rect 50820 36036 50848 36092
rect 50528 34524 50848 36036
rect 50528 34468 50556 34524
rect 50612 34468 50660 34524
rect 50716 34468 50764 34524
rect 50820 34468 50848 34524
rect 50528 32956 50848 34468
rect 50528 32900 50556 32956
rect 50612 32900 50660 32956
rect 50716 32900 50764 32956
rect 50820 32900 50848 32956
rect 50528 31388 50848 32900
rect 50528 31332 50556 31388
rect 50612 31332 50660 31388
rect 50716 31332 50764 31388
rect 50820 31332 50848 31388
rect 50528 29820 50848 31332
rect 50528 29764 50556 29820
rect 50612 29764 50660 29820
rect 50716 29764 50764 29820
rect 50820 29764 50848 29820
rect 50528 28252 50848 29764
rect 50528 28196 50556 28252
rect 50612 28196 50660 28252
rect 50716 28196 50764 28252
rect 50820 28196 50848 28252
rect 50528 26684 50848 28196
rect 50528 26628 50556 26684
rect 50612 26628 50660 26684
rect 50716 26628 50764 26684
rect 50820 26628 50848 26684
rect 50528 25116 50848 26628
rect 50528 25060 50556 25116
rect 50612 25060 50660 25116
rect 50716 25060 50764 25116
rect 50820 25060 50848 25116
rect 50528 23548 50848 25060
rect 50528 23492 50556 23548
rect 50612 23492 50660 23548
rect 50716 23492 50764 23548
rect 50820 23492 50848 23548
rect 50528 21980 50848 23492
rect 50528 21924 50556 21980
rect 50612 21924 50660 21980
rect 50716 21924 50764 21980
rect 50820 21924 50848 21980
rect 50528 20412 50848 21924
rect 50528 20356 50556 20412
rect 50612 20356 50660 20412
rect 50716 20356 50764 20412
rect 50820 20356 50848 20412
rect 50528 18844 50848 20356
rect 50528 18788 50556 18844
rect 50612 18788 50660 18844
rect 50716 18788 50764 18844
rect 50820 18788 50848 18844
rect 50528 17276 50848 18788
rect 50528 17220 50556 17276
rect 50612 17220 50660 17276
rect 50716 17220 50764 17276
rect 50820 17220 50848 17276
rect 50528 15708 50848 17220
rect 50528 15652 50556 15708
rect 50612 15652 50660 15708
rect 50716 15652 50764 15708
rect 50820 15652 50848 15708
rect 50528 14140 50848 15652
rect 50528 14084 50556 14140
rect 50612 14084 50660 14140
rect 50716 14084 50764 14140
rect 50820 14084 50848 14140
rect 50528 12572 50848 14084
rect 50528 12516 50556 12572
rect 50612 12516 50660 12572
rect 50716 12516 50764 12572
rect 50820 12516 50848 12572
rect 50528 11004 50848 12516
rect 50528 10948 50556 11004
rect 50612 10948 50660 11004
rect 50716 10948 50764 11004
rect 50820 10948 50848 11004
rect 50528 9436 50848 10948
rect 50528 9380 50556 9436
rect 50612 9380 50660 9436
rect 50716 9380 50764 9436
rect 50820 9380 50848 9436
rect 50528 7868 50848 9380
rect 50528 7812 50556 7868
rect 50612 7812 50660 7868
rect 50716 7812 50764 7868
rect 50820 7812 50848 7868
rect 50528 6300 50848 7812
rect 50528 6244 50556 6300
rect 50612 6244 50660 6300
rect 50716 6244 50764 6300
rect 50820 6244 50848 6300
rect 50528 4732 50848 6244
rect 50528 4676 50556 4732
rect 50612 4676 50660 4732
rect 50716 4676 50764 4732
rect 50820 4676 50848 4732
rect 50528 3164 50848 4676
rect 50528 3108 50556 3164
rect 50612 3108 50660 3164
rect 50716 3108 50764 3164
rect 50820 3108 50848 3164
rect 50528 3076 50848 3108
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _0563_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 25088 0 -1 50176
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__and4_1  _0564_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 36288 0 -1 53312
box -86 -86 1318 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_2  _0565_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 42224 0 1 51744
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_4  _0566_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 38192 0 1 51744
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_3  _0567_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform -1 0 38640 0 -1 31360
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _0568_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform -1 0 40096 0 -1 37632
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_3  _0569_
timestamp 1698175906
transform 1 0 32928 0 -1 34496
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _0570_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 38416 0 -1 37632
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_3  _0571_
timestamp 1698175906
transform -1 0 38640 0 -1 32928
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_3  _0572_
timestamp 1698175906
transform -1 0 39760 0 -1 34496
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__nand4_4  _0573_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 31920 0 1 32928
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _0574_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform -1 0 7280 0 1 48608
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _0575_
timestamp 1698175906
transform -1 0 6832 0 -1 48608
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _0576_
timestamp 1698175906
transform 1 0 7392 0 -1 50176
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _0577_
timestamp 1698175906
transform 1 0 8288 0 -1 50176
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _0578_
timestamp 1698175906
transform 1 0 3360 0 -1 48608
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _0579_
timestamp 1698175906
transform 1 0 8064 0 1 47040
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _0580_
timestamp 1698175906
transform 1 0 2016 0 1 47040
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  _0581_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 4368 0 -1 47040
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _0582_
timestamp 1698175906
transform 1 0 9520 0 -1 48608
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand4_2  _0583_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 10416 0 -1 48608
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_2  _0584_
timestamp 1698175906
transform -1 0 15456 0 -1 47040
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_3  _0585_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 24864 0 1 43904
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _0586_
timestamp 1698175906
transform 1 0 40768 0 -1 36064
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _0587_
timestamp 1698175906
transform -1 0 39984 0 -1 36064
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__inv_1  _0588_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 40096 0 -1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__buf_3  _0589_
timestamp 1698175906
transform -1 0 41104 0 1 36064
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_3  _0590_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 35728 0 1 32928
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _0591_
timestamp 1698175906
transform 1 0 40768 0 -1 32928
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _0592_
timestamp 1698175906
transform -1 0 34944 0 -1 37632
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor4_4  _0593_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 33152 0 -1 36064
box -86 -86 4230 870
use gf180mcu_fd_sc_mcu7t5v0__buf_3  _0594_
timestamp 1698175906
transform -1 0 31136 0 1 34496
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _0595_
timestamp 1698175906
transform 1 0 2800 0 -1 47040
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _0596_
timestamp 1698175906
transform 1 0 3360 0 -1 43904
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _0597_
timestamp 1698175906
transform 1 0 3808 0 1 47040
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _0598_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform -1 0 7392 0 -1 48608
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _0599_
timestamp 1698175906
transform 1 0 7952 0 1 45472
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_2  _0600_
timestamp 1698175906
transform -1 0 10192 0 1 40768
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__or2_1  _0601_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 6944 0 1 50176
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _0602_
timestamp 1698175906
transform -1 0 7952 0 1 45472
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_2  _0603_
timestamp 1698175906
transform -1 0 12320 0 1 43904
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__inv_2  _0604_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform -1 0 6720 0 -1 50176
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor4_4  _0605_
timestamp 1698175906
transform 1 0 8960 0 1 47040
box -86 -86 4230 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _0606_
timestamp 1698175906
transform 1 0 14112 0 -1 40768
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _0607_
timestamp 1698175906
transform -1 0 6944 0 1 47040
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  _0608_
timestamp 1698175906
transform -1 0 7392 0 -1 50176
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_3  _0609_
timestamp 1698175906
transform -1 0 7056 0 1 43904
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _0610_
timestamp 1698175906
transform 1 0 3808 0 1 45472
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor4_4  _0611_
timestamp 1698175906
transform -1 0 9184 0 -1 42336
box -86 -86 4230 870
use gf180mcu_fd_sc_mcu7t5v0__or4_1  _0612_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 13440 0 1 40768
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_2  _0613_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 3248 0 -1 47040
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _0614_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 6384 0 1 45472
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _0615_
timestamp 1698175906
transform -1 0 6384 0 1 37632
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _0616_
timestamp 1698175906
transform 1 0 13776 0 -1 39200
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_3  _0617_
timestamp 1698175906
transform 1 0 38416 0 1 36064
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__nor4_4  _0618_
timestamp 1698175906
transform 1 0 36848 0 1 34496
box -86 -86 4230 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _0619_
timestamp 1698175906
transform -1 0 12656 0 -1 34496
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _0620_
timestamp 1698175906
transform -1 0 12768 0 -1 29792
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_4  _0621_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform -1 0 39088 0 -1 36064
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  _0622_
timestamp 1698175906
transform -1 0 36176 0 1 29792
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _0623_
timestamp 1698175906
transform -1 0 35280 0 1 29792
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _0624_
timestamp 1698175906
transform -1 0 33488 0 1 36064
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _0625_
timestamp 1698175906
transform -1 0 32368 0 1 37632
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__or2_1  _0626_
timestamp 1698175906
transform 1 0 2912 0 1 47040
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _0627_
timestamp 1698175906
transform -1 0 5152 0 -1 43904
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__or2_2  _0628_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 11536 0 -1 40768
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _0629_
timestamp 1698175906
transform -1 0 11088 0 1 40768
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _0630_
timestamp 1698175906
transform 1 0 7168 0 1 47040
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _0631_
timestamp 1698175906
transform 1 0 3360 0 -1 42336
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand4_4  _0632_
timestamp 1698175906
transform 1 0 6272 0 1 39200
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _0633_
timestamp 1698175906
transform -1 0 33600 0 1 37632
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _0634_
timestamp 1698175906
transform -1 0 32480 0 1 36064
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand4_2  _0635_
timestamp 1698175906
transform -1 0 32704 0 -1 39200
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__oai32_2  _0636_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform -1 0 32144 0 1 39200
box -86 -86 2662 870
use gf180mcu_fd_sc_mcu7t5v0__aoi221_4  _0637_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform -1 0 19264 0 1 39200
box -86 -86 4566 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _0638_
timestamp 1698175906
transform 1 0 15008 0 1 43904
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_3  _0639_
timestamp 1698175906
transform -1 0 38416 0 1 36064
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__inv_1  _0640_
timestamp 1698175906
transform 1 0 36960 0 1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_3  _0641_
timestamp 1698175906
transform 1 0 38640 0 -1 32928
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__nor4_4  _0642_
timestamp 1698175906
transform 1 0 34160 0 -1 29792
box -86 -86 4230 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _0643_
timestamp 1698175906
transform -1 0 30800 0 -1 28224
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _0644_
timestamp 1698175906
transform 1 0 28000 0 1 28224
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _0645_
timestamp 1698175906
transform 1 0 21168 0 1 42336
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor4_4  _0646_
timestamp 1698175906
transform 1 0 37408 0 1 32928
box -86 -86 4230 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _0647_
timestamp 1698175906
transform -1 0 25984 0 -1 25088
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor4_4  _0648_
timestamp 1698175906
transform -1 0 40992 0 1 31360
box -86 -86 4230 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_3  _0649_
timestamp 1698175906
transform -1 0 31360 0 1 29792
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _0650_
timestamp 1698175906
transform 1 0 5152 0 -1 43904
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_4  _0651_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 5712 0 1 40768
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _0652_
timestamp 1698175906
transform -1 0 8064 0 -1 34496
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_2  _0653_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 23072 0 1 28224
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__nor4_2  _0654_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform -1 0 36624 0 1 34496
box -86 -86 2102 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _0655_
timestamp 1698175906
transform -1 0 31024 0 1 32928
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_4  _0656_
timestamp 1698175906
transform 1 0 34496 0 -1 34496
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _0657_
timestamp 1698175906
transform 1 0 27664 0 1 25088
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_4  _0658_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform -1 0 11536 0 -1 40768
box -86 -86 2102 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _0659_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform -1 0 28112 0 -1 29792
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_2  _0660_
timestamp 1698175906
transform -1 0 8624 0 1 42336
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _0661_
timestamp 1698175906
transform 1 0 22064 0 -1 39200
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_2  _0662_
timestamp 1698175906
transform -1 0 7840 0 -1 45472
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _0663_
timestamp 1698175906
transform 1 0 14112 0 1 43904
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _0664_
timestamp 1698175906
transform -1 0 30016 0 1 34496
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _0665_
timestamp 1698175906
transform 1 0 28560 0 -1 31360
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__and4_2  _0666_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 29008 0 1 28224
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_4  _0667_
timestamp 1698175906
transform 1 0 10192 0 1 45472
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _0668_
timestamp 1698175906
transform 1 0 14112 0 -1 32928
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_2  _0669_
timestamp 1698175906
transform 1 0 22400 0 1 29792
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_3  _0670_
timestamp 1698175906
transform 1 0 6384 0 1 34496
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__nor4_4  _0671_
timestamp 1698175906
transform 1 0 8624 0 1 42336
box -86 -86 4230 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _0672_
timestamp 1698175906
transform 1 0 9408 0 -1 34496
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_4  _0673_
timestamp 1698175906
transform -1 0 36400 0 1 36064
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _0674_
timestamp 1698175906
transform -1 0 25984 0 -1 31360
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_4  _0675_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform -1 0 28112 0 -1 32928
box -86 -86 3110 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _0676_
timestamp 1698175906
transform -1 0 30912 0 -1 34496
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _0677_
timestamp 1698175906
transform 1 0 11648 0 -1 37632
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _0678_
timestamp 1698175906
transform 1 0 7504 0 -1 28224
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _0679_
timestamp 1698175906
transform 1 0 20272 0 1 28224
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _0680_
timestamp 1698175906
transform -1 0 26320 0 1 26656
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _0681_
timestamp 1698175906
transform -1 0 24640 0 -1 29792
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__and4_1  _0682_
timestamp 1698175906
transform 1 0 24864 0 1 29792
box -86 -86 1318 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_4  _0683_
timestamp 1698175906
transform -1 0 28112 0 1 42336
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_3  _0684_
timestamp 1698175906
transform -1 0 10976 0 -1 28224
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__nor4_4  _0685_
timestamp 1698175906
transform 1 0 32928 0 -1 32928
box -86 -86 4230 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _0686_
timestamp 1698175906
transform 1 0 11984 0 1 26656
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _0687_
timestamp 1698175906
transform 1 0 7056 0 -1 43904
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _0688_
timestamp 1698175906
transform 1 0 7952 0 1 43904
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _0689_
timestamp 1698175906
transform 1 0 9520 0 1 48608
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand4_4  _0690_
timestamp 1698175906
transform 1 0 9632 0 -1 47040
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__oai31_2  _0691_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform -1 0 12992 0 -1 43904
box -86 -86 2214 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_4  _0692_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 11760 0 -1 28224
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_2  _0693_
timestamp 1698175906
transform -1 0 16128 0 1 47040
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _0694_
timestamp 1698175906
transform -1 0 16688 0 1 48608
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nor4_4  _0695_
timestamp 1698175906
transform -1 0 9184 0 -1 47040
box -86 -86 4230 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _0696_
timestamp 1698175906
transform 1 0 5488 0 1 36064
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor4_4  _0697_
timestamp 1698175906
transform -1 0 37072 0 -1 31360
box -86 -86 4230 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_3  _0698_
timestamp 1698175906
transform -1 0 24080 0 -1 32928
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__oai31_2  _0699_
timestamp 1698175906
transform -1 0 8736 0 1 36064
box -86 -86 2214 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_2  _0700_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform -1 0 16912 0 -1 40768
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__or3_1  _0701_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform -1 0 14560 0 -1 48608
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _0702_
timestamp 1698175906
transform -1 0 13888 0 -1 47040
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_4  _0703_
timestamp 1698175906
transform -1 0 34384 0 1 34496
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _0704_
timestamp 1698175906
transform -1 0 21728 0 -1 29792
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _0705_
timestamp 1698175906
transform -1 0 4480 0 -1 45472
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi211_2  _0706_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 6384 0 1 37632
box -86 -86 1990 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _0707_
timestamp 1698175906
transform -1 0 10752 0 -1 50176
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__or4_2  _0708_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform -1 0 38640 0 1 37632
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _0709_
timestamp 1698175906
transform -1 0 4032 0 -1 39200
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor4_2  _0710_
timestamp 1698175906
transform 1 0 5488 0 -1 39200
box -86 -86 2102 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _0711_
timestamp 1698175906
transform -1 0 4032 0 -1 34496
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _0712_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 6048 0 1 29792
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _0713_
timestamp 1698175906
transform -1 0 9184 0 -1 32928
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _0714_
timestamp 1698175906
transform -1 0 32256 0 1 29792
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _0715_
timestamp 1698175906
transform 1 0 6384 0 -1 43904
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _0716_
timestamp 1698175906
transform 1 0 7056 0 -1 25088
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _0717_
timestamp 1698175906
transform -1 0 12096 0 -1 26656
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _0718_
timestamp 1698175906
transform -1 0 12320 0 1 29792
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__and3_1  _0719_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 10640 0 1 34496
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__inv_1  _0720_
timestamp 1698175906
transform -1 0 20272 0 1 45472
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _0721_
timestamp 1698175906
transform -1 0 18368 0 1 42336
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor4_4  _0722_
timestamp 1698175906
transform 1 0 31920 0 1 31360
box -86 -86 4230 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _0723_
timestamp 1698175906
transform -1 0 23968 0 -1 39200
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _0724_
timestamp 1698175906
transform 1 0 22848 0 1 43904
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_2  _0725_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 17808 0 -1 48608
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nand4_4  _0726_
timestamp 1698175906
transform -1 0 20944 0 1 43904
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _0727_
timestamp 1698175906
transform -1 0 24976 0 1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _0728_
timestamp 1698175906
transform -1 0 24080 0 1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _0729_
timestamp 1698175906
transform 1 0 15568 0 1 26656
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _0730_
timestamp 1698175906
transform 1 0 13664 0 -1 36064
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _0731_
timestamp 1698175906
transform -1 0 29904 0 -1 28224
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _0732_
timestamp 1698175906
transform -1 0 6384 0 1 34496
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_2  _0733_
timestamp 1698175906
transform -1 0 16352 0 -1 34496
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__nand4_4  _0734_
timestamp 1698175906
transform 1 0 15120 0 1 34496
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _0735_
timestamp 1698175906
transform -1 0 3248 0 1 39200
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _0736_
timestamp 1698175906
transform -1 0 3584 0 1 31360
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor4_4  _0737_
timestamp 1698175906
transform 1 0 3472 0 -1 40768
box -86 -86 4230 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _0738_
timestamp 1698175906
transform -1 0 4480 0 1 31360
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _0739_
timestamp 1698175906
transform 1 0 33600 0 1 37632
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand4_4  _0740_
timestamp 1698175906
transform -1 0 35728 0 1 39200
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_2  _0741_
timestamp 1698175906
transform 1 0 11760 0 1 40768
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__nand4_4  _0742_
timestamp 1698175906
transform 1 0 33376 0 -1 39200
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__oai32_4  _0743_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 27888 0 -1 40768
box -86 -86 4902 870
use gf180mcu_fd_sc_mcu7t5v0__aoi221_4  _0744_
timestamp 1698175906
transform 1 0 2128 0 -1 29792
box -86 -86 4566 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _0745_
timestamp 1698175906
transform -1 0 12320 0 -1 36064
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _0746_
timestamp 1698175906
transform 1 0 5712 0 1 26656
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _0747_
timestamp 1698175906
transform -1 0 5264 0 1 29792
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nor4_2  _0748_
timestamp 1698175906
transform 1 0 3248 0 1 39200
box -86 -86 2102 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _0749_
timestamp 1698175906
transform -1 0 2912 0 -1 39200
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _0750_
timestamp 1698175906
transform 1 0 2352 0 1 37632
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__and3_1  _0751_
timestamp 1698175906
transform 1 0 4144 0 1 32928
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _0752_
timestamp 1698175906
transform -1 0 10640 0 1 34496
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_1  _0753_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 9408 0 -1 43904
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _0754_
timestamp 1698175906
transform 1 0 13328 0 1 42336
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _0755_
timestamp 1698175906
transform -1 0 12992 0 -1 26656
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_4  _0756_
timestamp 1698175906
transform 1 0 9968 0 -1 32928
box -86 -86 3110 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_3  _0757_
timestamp 1698175906
transform -1 0 14896 0 1 23520
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _0758_
timestamp 1698175906
transform -1 0 9296 0 1 25088
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _0759_
timestamp 1698175906
transform -1 0 14224 0 1 31360
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_4  _0760_
timestamp 1698175906
transform -1 0 12992 0 -1 31360
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__nand4_4  _0761_
timestamp 1698175906
transform -1 0 9408 0 1 32928
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__nor4_4  _0762_
timestamp 1698175906
transform 1 0 15456 0 1 40768
box -86 -86 4230 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _0763_
timestamp 1698175906
transform -1 0 19152 0 1 25088
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _0764_
timestamp 1698175906
transform -1 0 19376 0 -1 23520
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__aoi222_4  _0765_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 11760 0 -1 25088
box -86 -86 5350 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_3  _0766_
timestamp 1698175906
transform 1 0 21168 0 1 39200
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _0767_
timestamp 1698175906
transform 1 0 13776 0 -1 43904
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _0768_
timestamp 1698175906
transform -1 0 15792 0 1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_2  _0769_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform -1 0 22848 0 1 23520
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _0770_
timestamp 1698175906
transform 1 0 13664 0 -1 45472
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_2  _0771_
timestamp 1698175906
transform 1 0 19264 0 1 25088
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__nand4_4  _0772_
timestamp 1698175906
transform -1 0 21280 0 -1 25088
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _0773_
timestamp 1698175906
transform 1 0 7952 0 1 34496
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _0774_
timestamp 1698175906
transform 1 0 21952 0 -1 26656
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_2  _0775_
timestamp 1698175906
transform 1 0 20272 0 -1 36064
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _0776_
timestamp 1698175906
transform 1 0 5600 0 -1 36064
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_4  _0777_
timestamp 1698175906
transform 1 0 21504 0 1 34496
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _0778_
timestamp 1698175906
transform 1 0 7168 0 -1 26656
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi222_4  _0779_
timestamp 1698175906
transform -1 0 26880 0 1 25088
box -86 -86 5350 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_1  _0780_
timestamp 1698175906
transform -1 0 8400 0 -1 39200
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _0781_
timestamp 1698175906
transform -1 0 8064 0 -1 37632
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_2  _0782_
timestamp 1698175906
transform 1 0 30240 0 -1 37632
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__aoi222_4  _0783_
timestamp 1698175906
transform -1 0 27328 0 1 36064
box -86 -86 5350 870
use gf180mcu_fd_sc_mcu7t5v0__nand4_4  _0784_
timestamp 1698175906
transform -1 0 24864 0 -1 36064
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _0785_
timestamp 1698175906
transform 1 0 7504 0 -1 36064
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _0786_
timestamp 1698175906
transform 1 0 20048 0 1 34496
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _0787_
timestamp 1698175906
transform -1 0 31136 0 1 31360
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi222_2  _0788_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 19712 0 -1 34496
box -86 -86 2886 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _0789_
timestamp 1698175906
transform -1 0 20272 0 -1 36064
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _0790_
timestamp 1698175906
transform -1 0 13664 0 -1 31360
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _0791_
timestamp 1698175906
transform -1 0 29904 0 1 31360
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _0792_
timestamp 1698175906
transform 1 0 18256 0 -1 34496
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi222_4  _0793_
timestamp 1698175906
transform -1 0 24864 0 -1 37632
box -86 -86 5350 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_2  _0794_
timestamp 1698175906
transform 1 0 25088 0 -1 36064
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__nor4_4  _0795_
timestamp 1698175906
transform 1 0 23968 0 1 37632
box -86 -86 4230 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _0796_
timestamp 1698175906
transform 1 0 7840 0 -1 45472
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _0797_
timestamp 1698175906
transform 1 0 11648 0 -1 39200
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _0798_
timestamp 1698175906
transform -1 0 27888 0 -1 28224
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_2  _0799_
timestamp 1698175906
transform -1 0 25648 0 1 26656
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _0800_
timestamp 1698175906
transform -1 0 28000 0 -1 36064
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_2  _0801_
timestamp 1698175906
transform -1 0 26768 0 -1 37632
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__oai31_1  _0802_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform -1 0 8064 0 1 25088
box -86 -86 1318 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_2  _0803_
timestamp 1698175906
transform -1 0 9184 0 -1 40768
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _0804_
timestamp 1698175906
transform 1 0 9296 0 1 25088
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _0805_
timestamp 1698175906
transform -1 0 13104 0 1 25088
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_4  _0806_
timestamp 1698175906
transform 1 0 9520 0 -1 45472
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _0807_
timestamp 1698175906
transform 1 0 9184 0 1 45472
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_2  _0808_
timestamp 1698175906
transform -1 0 11648 0 1 39200
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _0809_
timestamp 1698175906
transform 1 0 11648 0 1 25088
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__and4_2  _0810_
timestamp 1698175906
transform 1 0 10192 0 1 25088
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _0811_
timestamp 1698175906
transform 1 0 23296 0 -1 43904
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__and4_1  _0812_
timestamp 1698175906
transform 1 0 25984 0 1 43904
box -86 -86 1318 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_4  _0813_
timestamp 1698175906
transform -1 0 28784 0 1 47040
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _0814_
timestamp 1698175906
transform 1 0 26320 0 -1 48608
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _0815_
timestamp 1698175906
transform 1 0 25424 0 -1 45472
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_2  _0816_
timestamp 1698175906
transform 1 0 23856 0 1 43904
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _0817_
timestamp 1698175906
transform 1 0 15792 0 1 50176
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__or3_1  _0818_
timestamp 1698175906
transform 1 0 13440 0 1 47040
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_2  _0819_
timestamp 1698175906
transform -1 0 26768 0 -1 34496
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_2  _0820_
timestamp 1698175906
transform -1 0 18928 0 -1 32928
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__oai211_1  _0821_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 15904 0 1 45472
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_2  _0822_
timestamp 1698175906
transform 1 0 18704 0 -1 45472
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _0823_
timestamp 1698175906
transform -1 0 17808 0 -1 48608
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _0824_
timestamp 1698175906
transform 1 0 17024 0 1 47040
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _0825_
timestamp 1698175906
transform -1 0 23072 0 1 31360
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_2  _0826_
timestamp 1698175906
transform -1 0 18704 0 1 32928
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_2  _0827_
timestamp 1698175906
transform -1 0 16128 0 1 37632
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__oai211_1  _0828_
timestamp 1698175906
transform 1 0 17248 0 -1 43904
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _0829_
timestamp 1698175906
transform -1 0 3360 0 1 32928
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _0830_
timestamp 1698175906
transform 1 0 2128 0 -1 36064
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _0831_
timestamp 1698175906
transform 1 0 3360 0 1 32928
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _0832_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 9744 0 -1 36064
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__aoi222_1  _0833_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 19376 0 1 31360
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _0834_
timestamp 1698175906
transform 1 0 12992 0 -1 32928
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _0835_
timestamp 1698175906
transform 1 0 14448 0 1 31360
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _0836_
timestamp 1698175906
transform 1 0 16016 0 -1 31360
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _0837_
timestamp 1698175906
transform 1 0 17360 0 -1 37632
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _0838_
timestamp 1698175906
transform 1 0 16464 0 -1 42336
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand4_1  _0839_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 17248 0 -1 31360
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__or4_1  _0840_
timestamp 1698175906
transform 1 0 16016 0 1 43904
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _0841_
timestamp 1698175906
transform -1 0 32480 0 -1 37632
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _0842_
timestamp 1698175906
transform -1 0 30240 0 -1 37632
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _0843_
timestamp 1698175906
transform 1 0 28224 0 1 36064
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai31_1  _0844_
timestamp 1698175906
transform -1 0 30800 0 1 37632
box -86 -86 1318 870
use gf180mcu_fd_sc_mcu7t5v0__nand4_4  _0845_
timestamp 1698175906
transform 1 0 10416 0 -1 42336
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _0846_
timestamp 1698175906
transform 1 0 12656 0 -1 40768
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_2  _0847_
timestamp 1698175906
transform 1 0 21504 0 -1 32928
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_4  _0848_
timestamp 1698175906
transform -1 0 24864 0 -1 25088
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__nand4_4  _0849_
timestamp 1698175906
transform 1 0 23520 0 1 31360
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _0850_
timestamp 1698175906
transform -1 0 12656 0 1 34496
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _0851_
timestamp 1698175906
transform -1 0 25760 0 -1 37632
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _0852_
timestamp 1698175906
transform 1 0 11536 0 1 37632
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _0853_
timestamp 1698175906
transform 1 0 12544 0 -1 39200
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand4_1  _0854_
timestamp 1698175906
transform -1 0 14336 0 1 37632
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__or4_1  _0855_
timestamp 1698175906
transform -1 0 26432 0 -1 39200
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__nor4_4  _0856_
timestamp 1698175906
transform 1 0 25984 0 -1 45472
box -86 -86 4230 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_4  _0857_
timestamp 1698175906
transform 1 0 26768 0 -1 48608
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _0858_
timestamp 1698175906
transform 1 0 24416 0 1 48608
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _0859_
timestamp 1698175906
transform -1 0 23632 0 1 32928
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_2  _0860_
timestamp 1698175906
transform -1 0 26544 0 1 34496
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _0861_
timestamp 1698175906
transform 1 0 27440 0 1 34496
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _0862_
timestamp 1698175906
transform -1 0 28448 0 1 32928
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _0863_
timestamp 1698175906
transform 1 0 28000 0 -1 36064
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_1  _0864_
timestamp 1698175906
transform -1 0 28672 0 1 39200
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _0865_
timestamp 1698175906
transform -1 0 3808 0 1 37632
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi222_4  _0866_
timestamp 1698175906
transform 1 0 1792 0 -1 32928
box -86 -86 5350 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _0867_
timestamp 1698175906
transform 1 0 5264 0 -1 34496
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _0868_
timestamp 1698175906
transform 1 0 18144 0 -1 37632
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _0869_
timestamp 1698175906
transform -1 0 19264 0 1 32928
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_2  _0870_
timestamp 1698175906
transform 1 0 12768 0 -1 34496
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _0871_
timestamp 1698175906
transform 1 0 2352 0 -1 37632
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _0872_
timestamp 1698175906
transform 1 0 16016 0 1 28224
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _0873_
timestamp 1698175906
transform -1 0 17808 0 -1 34496
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand4_1  _0874_
timestamp 1698175906
transform 1 0 16912 0 1 37632
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_4  _0875_
timestamp 1698175906
transform 1 0 17360 0 1 29792
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _0876_
timestamp 1698175906
transform 1 0 25760 0 1 28224
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _0877_
timestamp 1698175906
transform -1 0 18928 0 1 28224
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _0878_
timestamp 1698175906
transform -1 0 21840 0 -1 23520
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _0879_
timestamp 1698175906
transform -1 0 22624 0 1 28224
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _0880_
timestamp 1698175906
transform 1 0 18144 0 1 26656
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _0881_
timestamp 1698175906
transform -1 0 26096 0 -1 26656
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _0882_
timestamp 1698175906
transform -1 0 10304 0 1 37632
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _0883_
timestamp 1698175906
transform 1 0 17248 0 -1 26656
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__nand4_1  _0884_
timestamp 1698175906
transform 1 0 17584 0 -1 28224
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__nor4_1  _0885_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 18144 0 1 37632
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_2  _0886_
timestamp 1698175906
transform 1 0 9632 0 1 43904
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _0887_
timestamp 1698175906
transform 1 0 17696 0 -1 42336
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _0888_
timestamp 1698175906
transform -1 0 20160 0 1 40768
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _0889_
timestamp 1698175906
transform 1 0 17920 0 1 48608
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_1  _0890_
timestamp 1698175906
transform 1 0 17920 0 1 47040
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _0891_
timestamp 1698175906
transform -1 0 18480 0 1 36064
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_1  _0892_
timestamp 1698175906
transform 1 0 18256 0 -1 42336
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__and4_1  _0893_
timestamp 1698175906
transform 1 0 18368 0 -1 40768
box -86 -86 1318 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_2  _0894_
timestamp 1698175906
transform -1 0 24640 0 1 45472
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__nand4_2  _0895_
timestamp 1698175906
transform -1 0 29904 0 -1 29792
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _0896_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 26320 0 -1 28224
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _0897_
timestamp 1698175906
transform -1 0 28672 0 -1 32928
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_2  _0898_
timestamp 1698175906
transform -1 0 19264 0 1 31360
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _0899_
timestamp 1698175906
transform -1 0 28224 0 -1 31360
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_2  _0900_
timestamp 1698175906
transform 1 0 27104 0 1 31360
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__or4_1  _0901_
timestamp 1698175906
transform -1 0 28112 0 -1 37632
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _0902_
timestamp 1698175906
transform -1 0 6272 0 -1 26656
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__or2_1  _0903_
timestamp 1698175906
transform 1 0 8176 0 -1 34496
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _0904_
timestamp 1698175906
transform 1 0 13328 0 1 25088
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi222_4  _0905_
timestamp 1698175906
transform 1 0 7840 0 1 31360
box -86 -86 5350 870
use gf180mcu_fd_sc_mcu7t5v0__oai31_1  _0906_
timestamp 1698175906
transform -1 0 14112 0 -1 29792
box -86 -86 1318 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _0907_
timestamp 1698175906
transform 1 0 14560 0 1 28224
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _0908_
timestamp 1698175906
transform 1 0 13776 0 -1 31360
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__and3_1  _0909_
timestamp 1698175906
transform 1 0 14224 0 -1 29792
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nand4_4  _0910_
timestamp 1698175906
transform 1 0 23184 0 1 40768
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _0911_
timestamp 1698175906
transform 1 0 13776 0 1 45472
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _0912_
timestamp 1698175906
transform 1 0 21392 0 -1 48608
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _0913_
timestamp 1698175906
transform 1 0 22736 0 1 48608
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _0914_
timestamp 1698175906
transform 1 0 23744 0 -1 48608
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nor4_4  _0915_
timestamp 1698175906
transform 1 0 24640 0 1 45472
box -86 -86 4230 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_4  _0916_
timestamp 1698175906
transform -1 0 28448 0 1 48608
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _0917_
timestamp 1698175906
transform 1 0 27440 0 -1 50176
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _0918_
timestamp 1698175906
transform 1 0 24416 0 -1 43904
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _0919_
timestamp 1698175906
transform 1 0 23744 0 1 42336
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nor4_4  _0920_
timestamp 1698175906
transform 1 0 26432 0 -1 43904
box -86 -86 4230 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _0921_
timestamp 1698175906
transform 1 0 24304 0 1 42336
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _0922_
timestamp 1698175906
transform 1 0 25088 0 -1 28224
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _0923_
timestamp 1698175906
transform 1 0 18368 0 -1 31360
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _0924_
timestamp 1698175906
transform 1 0 25984 0 -1 31360
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _0925_
timestamp 1698175906
transform 1 0 24080 0 -1 31360
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_1  _0926_
timestamp 1698175906
transform -1 0 25984 0 -1 40768
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_2  _0927_
timestamp 1698175906
transform 1 0 23408 0 1 29792
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _0928_
timestamp 1698175906
transform -1 0 10864 0 -1 34496
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _0929_
timestamp 1698175906
transform -1 0 9184 0 -1 28224
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _0930_
timestamp 1698175906
transform -1 0 11536 0 1 28224
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__nand4_2  _0931_
timestamp 1698175906
transform -1 0 11200 0 -1 29792
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_2  _0932_
timestamp 1698175906
transform -1 0 8960 0 -1 29792
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_2  _0933_
timestamp 1698175906
transform 1 0 1904 0 -1 31360
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__nand4_4  _0934_
timestamp 1698175906
transform 1 0 3696 0 -1 31360
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _0935_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 2240 0 1 40768
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _0936_
timestamp 1698175906
transform 1 0 2912 0 -1 45472
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _0937_
timestamp 1698175906
transform 1 0 14224 0 1 25088
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _0938_
timestamp 1698175906
transform -1 0 21840 0 -1 26656
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _0939_
timestamp 1698175906
transform 1 0 8960 0 1 26656
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _0940_
timestamp 1698175906
transform 1 0 9408 0 -1 26656
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _0941_
timestamp 1698175906
transform -1 0 5712 0 -1 28224
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__nand4_2  _0942_
timestamp 1698175906
transform 1 0 5712 0 -1 28224
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__nor4_4  _0943_
timestamp 1698175906
transform 1 0 6384 0 1 28224
box -86 -86 4230 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _0944_
timestamp 1698175906
transform 1 0 17248 0 -1 40768
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _0945_
timestamp 1698175906
transform -1 0 21728 0 1 28224
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand4_2  _0946_
timestamp 1698175906
transform 1 0 22512 0 -1 34496
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _0947_
timestamp 1698175906
transform 1 0 18032 0 1 50176
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _0948_
timestamp 1698175906
transform 1 0 18592 0 1 48608
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi211_1  _0949_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform -1 0 22736 0 1 48608
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__and4_1  _0950_
timestamp 1698175906
transform 1 0 25088 0 -1 43904
box -86 -86 1318 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_4  _0951_
timestamp 1698175906
transform 1 0 29008 0 1 47040
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__inv_1  _0952_
timestamp 1698175906
transform -1 0 38864 0 1 45472
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__buf_3  _0953_
timestamp 1698175906
transform 1 0 27664 0 1 43904
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__and3_1  _0954_
timestamp 1698175906
transform 1 0 21168 0 1 43904
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nand4_1  _0955_
timestamp 1698175906
transform 1 0 20048 0 -1 42336
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__aoi221_1  _0956_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 21504 0 -1 45472
box -86 -86 1318 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_2  _0957_
timestamp 1698175906
transform 1 0 18592 0 -1 28224
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__nand4_1  _0958_
timestamp 1698175906
transform -1 0 19712 0 1 34496
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _0959_
timestamp 1698175906
transform 1 0 15232 0 -1 26656
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__nand4_2  _0960_
timestamp 1698175906
transform 1 0 15680 0 1 31360
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _0961_
timestamp 1698175906
transform -1 0 4368 0 -1 28224
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _0962_
timestamp 1698175906
transform 1 0 2352 0 -1 45472
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _0963_
timestamp 1698175906
transform 1 0 2128 0 1 34496
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _0964_
timestamp 1698175906
transform 1 0 3136 0 -1 36064
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__nor4_2  _0965_
timestamp 1698175906
transform 1 0 17472 0 -1 36064
box -86 -86 2102 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _0966_
timestamp 1698175906
transform 1 0 22736 0 -1 45472
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__and3_1  _0967_
timestamp 1698175906
transform -1 0 28560 0 -1 34496
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nand4_4  _0968_
timestamp 1698175906
transform -1 0 27216 0 1 32928
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__or2_1  _0969_
timestamp 1698175906
transform 1 0 25984 0 -1 40768
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor4_4  _0970_
timestamp 1698175906
transform -1 0 31808 0 -1 42336
box -86 -86 4230 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_4  _0971_
timestamp 1698175906
transform 1 0 29008 0 1 45472
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__inv_1  _0972_
timestamp 1698175906
transform -1 0 41216 0 -1 42336
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _0973_
timestamp 1698175906
transform 1 0 28112 0 1 37632
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _0974_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 26544 0 1 34496
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _0975_
timestamp 1698175906
transform 1 0 19712 0 1 47040
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _0976_
timestamp 1698175906
transform -1 0 20944 0 1 36064
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__and4_1  _0977_
timestamp 1698175906
transform 1 0 19488 0 1 37632
box -86 -86 1318 870
use gf180mcu_fd_sc_mcu7t5v0__and4_1  _0978_
timestamp 1698175906
transform 1 0 20832 0 -1 39200
box -86 -86 1318 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _0979_
timestamp 1698175906
transform -1 0 11536 0 1 37632
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__aoi222_2  _0980_
timestamp 1698175906
transform 1 0 7392 0 1 29792
box -86 -86 2886 870
use gf180mcu_fd_sc_mcu7t5v0__aoi222_2  _0981_
timestamp 1698175906
transform 1 0 1792 0 1 36064
box -86 -86 2886 870
use gf180mcu_fd_sc_mcu7t5v0__and4_1  _0982_
timestamp 1698175906
transform 1 0 9408 0 -1 37632
box -86 -86 1318 870
use gf180mcu_fd_sc_mcu7t5v0__and4_1  _0983_
timestamp 1698175906
transform 1 0 26432 0 -1 39200
box -86 -86 1318 870
use gf180mcu_fd_sc_mcu7t5v0__and3_1  _0984_
timestamp 1698175906
transform 1 0 19824 0 1 23520
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _0985_
timestamp 1698175906
transform -1 0 15568 0 1 26656
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _0986_
timestamp 1698175906
transform 1 0 16464 0 -1 28224
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__and3_1  _0987_
timestamp 1698175906
transform 1 0 15344 0 -1 28224
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_2  _0988_
timestamp 1698175906
transform -1 0 21728 0 -1 28224
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_2  _0989_
timestamp 1698175906
transform -1 0 18480 0 1 25088
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _0990_
timestamp 1698175906
transform 1 0 15680 0 -1 23520
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_2  _0991_
timestamp 1698175906
transform 1 0 15008 0 1 25088
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__nand4_4  _0992_
timestamp 1698175906
transform 1 0 16240 0 1 23520
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _0993_
timestamp 1698175906
transform 1 0 22624 0 -1 48608
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _0994_
timestamp 1698175906
transform 1 0 23184 0 -1 48608
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nor4_4  _0995_
timestamp 1698175906
transform 1 0 23184 0 1 39200
box -86 -86 4230 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_4  _0996_
timestamp 1698175906
transform 1 0 30912 0 1 40768
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _0997_
timestamp 1698175906
transform -1 0 38864 0 1 42336
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__oai211_2  _0998_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform -1 0 28784 0 1 40768
box -86 -86 2102 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_2  _0999_
timestamp 1698175906
transform 1 0 29008 0 1 43904
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1000_
timestamp 1698175906
transform 1 0 20384 0 1 40768
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1001_
timestamp 1698175906
transform 1 0 18928 0 -1 37632
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai31_1  _1002_
timestamp 1698175906
transform 1 0 19936 0 -1 31360
box -86 -86 1318 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _1003_
timestamp 1698175906
transform -1 0 20608 0 -1 29792
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__nand4_1  _1004_
timestamp 1698175906
transform 1 0 21168 0 1 29792
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__nor4_1  _1005_
timestamp 1698175906
transform 1 0 21168 0 1 40768
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_2  _1006_
timestamp 1698175906
transform 1 0 13328 0 1 34496
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _1007_
timestamp 1698175906
transform 1 0 2128 0 -1 42336
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _1008_
timestamp 1698175906
transform 1 0 3136 0 1 28224
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__and3_1  _1009_
timestamp 1698175906
transform -1 0 9184 0 -1 37632
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__and4_1  _1010_
timestamp 1698175906
transform 1 0 3808 0 1 37632
box -86 -86 1318 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1011_
timestamp 1698175906
transform 1 0 19824 0 -1 47040
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__or4_1  _1012_
timestamp 1698175906
transform 1 0 20160 0 -1 45472
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__aoi222_1  _1013_
timestamp 1698175906
transform 1 0 21168 0 1 45472
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__and4_1  _1014_
timestamp 1698175906
transform 1 0 21728 0 -1 42336
box -86 -86 1318 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_4  _1015_
timestamp 1698175906
transform 1 0 30688 0 1 42336
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1016_
timestamp 1698175906
transform -1 0 37744 0 1 43904
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__or3_1  _1017_
timestamp 1698175906
transform 1 0 29008 0 1 40768
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_2  _1018_
timestamp 1698175906
transform -1 0 30688 0 1 42336
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _1019_
timestamp 1698175906
transform -1 0 19600 0 1 47040
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1020_
timestamp 1698175906
transform -1 0 20720 0 1 48608
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_2  _1021_
timestamp 1698175906
transform -1 0 20384 0 -1 48608
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1022_
timestamp 1698175906
transform 1 0 12432 0 1 29792
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _1023_
timestamp 1698175906
transform -1 0 14448 0 1 36064
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1024_
timestamp 1698175906
transform 1 0 14560 0 -1 36064
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _1025_
timestamp 1698175906
transform 1 0 15904 0 -1 37632
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__nand4_1  _1026_
timestamp 1698175906
transform 1 0 14672 0 -1 39200
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__or3_1  _1027_
timestamp 1698175906
transform 1 0 14784 0 -1 37632
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _1028_
timestamp 1698175906
transform 1 0 2128 0 -1 43904
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _1029_
timestamp 1698175906
transform -1 0 3136 0 1 28224
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1030_
timestamp 1698175906
transform 1 0 2576 0 1 42336
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nor4_4  _1031_
timestamp 1698175906
transform 1 0 18480 0 -1 43904
box -86 -86 4230 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_4  _1032_
timestamp 1698175906
transform 1 0 30464 0 1 43904
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__inv_1  _1033_
timestamp 1698175906
transform -1 0 23184 0 1 54880
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1034_
timestamp 1698175906
transform -1 0 10416 0 -1 53312
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1035_
timestamp 1698175906
transform 1 0 11648 0 1 54880
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_2  _1036_
timestamp 1698175906
transform 1 0 12992 0 -1 54880
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1037_
timestamp 1698175906
transform -1 0 12544 0 -1 53312
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1038_
timestamp 1698175906
transform 1 0 12656 0 -1 50176
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1039_
timestamp 1698175906
transform 1 0 11760 0 -1 50176
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi211_1  _1040_
timestamp 1698175906
transform 1 0 10528 0 -1 51744
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__inv_1  _1041_
timestamp 1698175906
transform -1 0 25536 0 1 54880
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1042_
timestamp 1698175906
transform 1 0 11088 0 -1 50176
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi211_1  _1043_
timestamp 1698175906
transform 1 0 9856 0 1 51744
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__inv_1  _1044_
timestamp 1698175906
transform -1 0 27888 0 1 54880
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1045_
timestamp 1698175906
transform 1 0 10976 0 1 48608
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi211_1  _1046_
timestamp 1698175906
transform 1 0 10416 0 -1 53312
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__inv_1  _1047_
timestamp 1698175906
transform -1 0 29904 0 -1 53312
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1048_
timestamp 1698175906
transform 1 0 31584 0 -1 43904
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1049_
timestamp 1698175906
transform 1 0 12992 0 -1 43904
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi211_1  _1050_
timestamp 1698175906
transform 1 0 10976 0 1 51744
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  _1051_
timestamp 1698175906
transform -1 0 32928 0 1 54880
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1052_
timestamp 1698175906
transform 1 0 32928 0 -1 43904
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1053_
timestamp 1698175906
transform -1 0 35392 0 1 50176
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1054_
timestamp 1698175906
transform 1 0 35728 0 1 40768
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi211_1  _1055_
timestamp 1698175906
transform 1 0 34832 0 -1 42336
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  _1056_
timestamp 1698175906
transform -1 0 34944 0 -1 54880
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1057_
timestamp 1698175906
transform 1 0 34160 0 -1 40768
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi211_1  _1058_
timestamp 1698175906
transform 1 0 34608 0 1 40768
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  _1059_
timestamp 1698175906
transform 1 0 36848 0 1 54880
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1060_
timestamp 1698175906
transform 1 0 34160 0 -1 42336
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi211_1  _1061_
timestamp 1698175906
transform 1 0 34832 0 -1 40768
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  _1062_
timestamp 1698175906
transform -1 0 39424 0 1 54880
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1063_
timestamp 1698175906
transform 1 0 33040 0 -1 45472
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi211_1  _1064_
timestamp 1698175906
transform -1 0 35168 0 1 43904
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_2  _1065_
timestamp 1698175906
transform 1 0 14784 0 -1 48608
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1066_
timestamp 1698175906
transform 1 0 21952 0 1 50176
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1067_
timestamp 1698175906
transform 1 0 24304 0 1 50176
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1068_
timestamp 1698175906
transform 1 0 12320 0 -1 54880
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1069_
timestamp 1698175906
transform -1 0 27216 0 -1 53312
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1070_
timestamp 1698175906
transform 1 0 23408 0 1 50176
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1071_
timestamp 1698175906
transform 1 0 22288 0 -1 53312
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1072_
timestamp 1698175906
transform 1 0 26096 0 1 53312
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1073_
timestamp 1698175906
transform 1 0 24528 0 1 53312
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1074_
timestamp 1698175906
transform 1 0 23408 0 1 53312
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1075_
timestamp 1698175906
transform 1 0 22176 0 1 53312
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1076_
timestamp 1698175906
transform -1 0 26320 0 -1 53312
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1077_
timestamp 1698175906
transform 1 0 26208 0 1 50176
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1078_
timestamp 1698175906
transform 1 0 37968 0 1 47040
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1079_
timestamp 1698175906
transform 1 0 38976 0 -1 47040
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1080_
timestamp 1698175906
transform 1 0 39088 0 -1 48608
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1081_
timestamp 1698175906
transform 1 0 38864 0 1 47040
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1082_
timestamp 1698175906
transform -1 0 41664 0 -1 47040
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1083_
timestamp 1698175906
transform 1 0 40992 0 -1 43904
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1084_
timestamp 1698175906
transform 1 0 40096 0 1 42336
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1085_
timestamp 1698175906
transform 1 0 38864 0 1 42336
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1086_
timestamp 1698175906
transform -1 0 39648 0 1 43904
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1087_
timestamp 1698175906
transform -1 0 40544 0 -1 45472
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1088_
timestamp 1698175906
transform -1 0 42112 0 1 45472
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1089_
timestamp 1698175906
transform 1 0 29008 0 -1 54880
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1090_
timestamp 1698175906
transform 1 0 32816 0 1 53312
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1091_
timestamp 1698175906
transform -1 0 38752 0 1 54880
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1092_
timestamp 1698175906
transform -1 0 32256 0 -1 54880
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi211_1  _1093_
timestamp 1698175906
transform 1 0 29680 0 -1 54880
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1094_
timestamp 1698175906
transform -1 0 32480 0 -1 53312
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi211_1  _1095_
timestamp 1698175906
transform 1 0 29904 0 -1 53312
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1096_
timestamp 1698175906
transform -1 0 36848 0 -1 54880
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi211_1  _1097_
timestamp 1698175906
transform 1 0 33040 0 -1 54880
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1098_
timestamp 1698175906
transform -1 0 38640 0 1 53312
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1099_
timestamp 1698175906
transform 1 0 37520 0 -1 53312
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi211_1  _1100_
timestamp 1698175906
transform 1 0 33040 0 -1 53312
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1101_
timestamp 1698175906
transform 1 0 38416 0 -1 54880
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1102_
timestamp 1698175906
transform 1 0 38640 0 1 53312
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1103_
timestamp 1698175906
transform -1 0 40432 0 -1 51744
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi211_1  _1104_
timestamp 1698175906
transform 1 0 38640 0 -1 51744
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1105_
timestamp 1698175906
transform -1 0 42672 0 1 53312
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi211_1  _1106_
timestamp 1698175906
transform 1 0 41104 0 1 51744
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1107_
timestamp 1698175906
transform -1 0 42672 0 -1 51744
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi211_1  _1108_
timestamp 1698175906
transform 1 0 40880 0 -1 51744
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1109_
timestamp 1698175906
transform 1 0 40768 0 1 53312
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi211_1  _1110_
timestamp 1698175906
transform -1 0 41888 0 -1 54880
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_2  _1111_
timestamp 1698175906
transform 1 0 15008 0 1 48608
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1112_
timestamp 1698175906
transform -1 0 17024 0 -1 51744
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1113_
timestamp 1698175906
transform -1 0 17920 0 -1 51744
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1114_
timestamp 1698175906
transform 1 0 16240 0 1 53312
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1115_
timestamp 1698175906
transform 1 0 15568 0 -1 54880
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1116_
timestamp 1698175906
transform 1 0 14560 0 -1 54880
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1117_
timestamp 1698175906
transform 1 0 15456 0 1 51744
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1118_
timestamp 1698175906
transform 1 0 14448 0 1 51744
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1119_
timestamp 1698175906
transform 1 0 18144 0 -1 54880
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1120_
timestamp 1698175906
transform 1 0 17248 0 -1 54880
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1121_
timestamp 1698175906
transform 1 0 18032 0 -1 51744
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1122_
timestamp 1698175906
transform 1 0 17920 0 -1 53312
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1123_
timestamp 1698175906
transform 1 0 30352 0 -1 48608
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1124_
timestamp 1698175906
transform 1 0 30240 0 1 50176
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1125_
timestamp 1698175906
transform 1 0 33040 0 1 47040
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1126_
timestamp 1698175906
transform 1 0 32592 0 1 45472
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1127_
timestamp 1698175906
transform -1 0 33824 0 -1 47040
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1128_
timestamp 1698175906
transform -1 0 34608 0 1 47040
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1129_
timestamp 1698175906
transform -1 0 35168 0 -1 50176
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1130_
timestamp 1698175906
transform -1 0 35056 0 1 45472
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1131_
timestamp 1698175906
transform -1 0 35504 0 1 47040
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1132_
timestamp 1698175906
transform 1 0 32928 0 -1 50176
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1133_
timestamp 1698175906
transform 1 0 31024 0 -1 48608
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1134_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform -1 0 4816 0 -1 50176
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1135_
timestamp 1698175906
transform -1 0 4816 0 1 50176
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1136_
timestamp 1698175906
transform -1 0 8960 0 -1 53312
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1137_
timestamp 1698175906
transform 1 0 4144 0 -1 51744
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1138_
timestamp 1698175906
transform 1 0 36848 0 -1 40768
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_2  _1139_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 34944 0 -1 37632
box -86 -86 3558 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1140_
timestamp 1698175906
transform 1 0 37296 0 -1 39200
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1141_
timestamp 1698175906
transform 1 0 33712 0 -1 43904
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1142_
timestamp 1698175906
transform 1 0 20832 0 -1 51744
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1143_
timestamp 1698175906
transform 1 0 25088 0 -1 54880
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1144_
timestamp 1698175906
transform 1 0 20832 0 -1 54880
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1145_
timestamp 1698175906
transform 1 0 25200 0 -1 51744
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1146_
timestamp 1698175906
transform -1 0 43008 0 1 47040
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1147_
timestamp 1698175906
transform 1 0 40992 0 1 42336
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1148_
timestamp 1698175906
transform -1 0 40320 0 -1 43904
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1149_
timestamp 1698175906
transform 1 0 41440 0 -1 45472
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1150_
timestamp 1698175906
transform 1 0 29008 0 1 54880
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1151_
timestamp 1698175906
transform 1 0 29232 0 1 51744
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1152_
timestamp 1698175906
transform 1 0 33376 0 1 54880
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1153_
timestamp 1698175906
transform 1 0 33264 0 1 51744
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1154_
timestamp 1698175906
transform 1 0 36960 0 1 50176
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1155_
timestamp 1698175906
transform 1 0 41776 0 -1 53312
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1156_
timestamp 1698175906
transform 1 0 41104 0 1 50176
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1157_
timestamp 1698175906
transform 1 0 40096 0 1 54880
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1158_
timestamp 1698175906
transform 1 0 13328 0 1 54880
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1159_
timestamp 1698175906
transform 1 0 12992 0 -1 51744
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1160_
timestamp 1698175906
transform 1 0 17472 0 1 54880
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1161_
timestamp 1698175906
transform -1 0 20944 0 1 51744
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1162_
timestamp 1698175906
transform -1 0 32704 0 1 48608
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1163_
timestamp 1698175906
transform -1 0 36624 0 1 48608
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1164_
timestamp 1698175906
transform -1 0 37632 0 -1 47040
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1165_
timestamp 1698175906
transform -1 0 32368 0 -1 50176
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0567__I $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform -1 0 37296 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0584__A1
timestamp 1698175906
transform 1 0 16128 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0584__A2
timestamp 1698175906
transform 1 0 15680 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0585__I
timestamp 1698175906
transform 1 0 24640 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0586__I
timestamp 1698175906
transform 1 0 40320 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0612__A3
timestamp 1698175906
transform 1 0 15008 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0619__I
timestamp 1698175906
transform 1 0 12880 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0622__I
timestamp 1698175906
transform -1 0 36624 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0636__A3
timestamp 1698175906
transform -1 0 29568 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0636__B1
timestamp 1698175906
transform -1 0 29344 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0637__A1
timestamp 1698175906
transform -1 0 20160 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0637__B1
timestamp 1698175906
transform -1 0 14784 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0637__B2
timestamp 1698175906
transform 1 0 14112 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0644__A1
timestamp 1698175906
transform 1 0 27328 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0644__A2
timestamp 1698175906
transform -1 0 28000 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0647__I
timestamp 1698175906
transform 1 0 26208 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0653__A1
timestamp 1698175906
transform 1 0 22848 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0653__B1
timestamp 1698175906
transform 1 0 25088 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0653__B2
timestamp 1698175906
transform 1 0 22624 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0657__I
timestamp 1698175906
transform 1 0 29232 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0659__A1
timestamp 1698175906
transform -1 0 27216 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0659__A2
timestamp 1698175906
transform 1 0 29232 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0659__B
timestamp 1698175906
transform 1 0 26544 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0665__A2
timestamp 1698175906
transform 1 0 28336 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0668__I
timestamp 1698175906
transform 1 0 13888 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0669__A1
timestamp 1698175906
transform -1 0 23632 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0674__I
timestamp 1698175906
transform 1 0 26320 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0675__A1
timestamp 1698175906
transform 1 0 24640 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0675__A2
timestamp 1698175906
transform -1 0 23520 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0677__I
timestamp 1698175906
transform 1 0 12544 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0679__A1
timestamp 1698175906
transform 1 0 20048 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0680__I
timestamp 1698175906
transform 1 0 26544 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0681__A1
timestamp 1698175906
transform 1 0 23856 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0683__A2
timestamp 1698175906
transform 1 0 28336 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0686__I
timestamp 1698175906
transform 1 0 13552 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0692__B2
timestamp 1698175906
transform 1 0 14448 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0693__A1
timestamp 1698175906
transform 1 0 16800 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0693__A2
timestamp 1698175906
transform 1 0 16352 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0699__B
timestamp 1698175906
transform 1 0 8960 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0700__A3
timestamp 1698175906
transform -1 0 15456 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0701__A1
timestamp 1698175906
transform 1 0 16576 0 -1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0701__A2
timestamp 1698175906
transform 1 0 16128 0 -1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0704__I
timestamp 1698175906
transform 1 0 21952 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0706__A2
timestamp 1698175906
transform -1 0 6384 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0708__A1
timestamp 1698175906
transform 1 0 36400 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0709__I
timestamp 1698175906
transform 1 0 4256 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0716__I
timestamp 1698175906
transform -1 0 7056 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0718__A2
timestamp 1698175906
transform -1 0 11872 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0718__B1
timestamp 1698175906
transform -1 0 11312 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0719__A1
timestamp 1698175906
transform 1 0 12544 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0723__I
timestamp 1698175906
transform -1 0 24192 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0726__A3
timestamp 1698175906
transform 1 0 20720 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0727__I
timestamp 1698175906
transform -1 0 25536 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0729__A2
timestamp 1698175906
transform -1 0 14784 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0733__A2
timestamp 1698175906
transform -1 0 16800 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0733__B1
timestamp 1698175906
transform 1 0 14112 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0733__B2
timestamp 1698175906
transform 1 0 16352 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0735__A1
timestamp 1698175906
transform -1 0 3472 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0737__A4
timestamp 1698175906
transform 1 0 6048 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0743__A3
timestamp 1698175906
transform 1 0 27552 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0743__B2
timestamp 1698175906
transform -1 0 27440 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0744__A1
timestamp 1698175906
transform 1 0 6160 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0744__C
timestamp 1698175906
transform 1 0 5824 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0745__A2
timestamp 1698175906
transform 1 0 12992 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0747__A1
timestamp 1698175906
transform -1 0 4704 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0747__A2
timestamp 1698175906
transform -1 0 4256 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0748__A3
timestamp 1698175906
transform 1 0 5264 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0752__I
timestamp 1698175906
transform 1 0 10752 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0755__I
timestamp 1698175906
transform 1 0 13216 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0756__A2
timestamp 1698175906
transform -1 0 13104 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0756__B
timestamp 1698175906
transform 1 0 12432 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0759__I
timestamp 1698175906
transform 1 0 15232 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0761__A3
timestamp 1698175906
transform 1 0 9632 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0763__I
timestamp 1698175906
transform 1 0 16800 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0765__A1
timestamp 1698175906
transform -1 0 11760 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0765__A2
timestamp 1698175906
transform -1 0 17696 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0768__I
timestamp 1698175906
transform -1 0 15232 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0769__A1
timestamp 1698175906
transform -1 0 23072 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0769__A2
timestamp 1698175906
transform -1 0 21168 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0771__A1
timestamp 1698175906
transform 1 0 19040 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0771__A2
timestamp 1698175906
transform -1 0 17696 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0771__B
timestamp 1698175906
transform 1 0 20272 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0774__I
timestamp 1698175906
transform 1 0 23072 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0777__A1
timestamp 1698175906
transform 1 0 21840 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0777__A2
timestamp 1698175906
transform 1 0 29680 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0777__B2
timestamp 1698175906
transform -1 0 21616 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0778__I
timestamp 1698175906
transform 1 0 6944 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0779__A1
timestamp 1698175906
transform -1 0 21616 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0779__B2
timestamp 1698175906
transform 1 0 19824 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0779__C1
timestamp 1698175906
transform 1 0 27104 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0779__C2
timestamp 1698175906
transform 1 0 20720 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0780__A3
timestamp 1698175906
transform 1 0 8624 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0783__A1
timestamp 1698175906
transform 1 0 29680 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0783__A2
timestamp 1698175906
transform 1 0 21504 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0783__B1
timestamp 1698175906
transform 1 0 19264 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0783__B2
timestamp 1698175906
transform -1 0 28560 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0783__C2
timestamp 1698175906
transform -1 0 19936 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0786__A1
timestamp 1698175906
transform 1 0 19824 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0786__A2
timestamp 1698175906
transform -1 0 20384 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0786__B
timestamp 1698175906
transform -1 0 19040 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0788__B1
timestamp 1698175906
transform 1 0 18032 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0788__B2
timestamp 1698175906
transform 1 0 19488 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0788__C1
timestamp 1698175906
transform 1 0 20272 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0788__C2
timestamp 1698175906
transform 1 0 19488 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0793__A1
timestamp 1698175906
transform 1 0 19376 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0793__A2
timestamp 1698175906
transform -1 0 22624 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0793__B1
timestamp 1698175906
transform 1 0 24192 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0793__C1
timestamp 1698175906
transform -1 0 19152 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0793__C2
timestamp 1698175906
transform -1 0 23520 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0795__A1
timestamp 1698175906
transform 1 0 21952 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0798__I
timestamp 1698175906
transform -1 0 27216 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0799__A2
timestamp 1698175906
transform 1 0 23744 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0800__I
timestamp 1698175906
transform 1 0 28784 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0801__A1
timestamp 1698175906
transform 1 0 24640 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0802__B
timestamp 1698175906
transform -1 0 8400 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0805__A2
timestamp 1698175906
transform -1 0 13104 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0809__A1
timestamp 1698175906
transform -1 0 11312 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0809__B
timestamp 1698175906
transform -1 0 11760 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0811__I
timestamp 1698175906
transform 1 0 22624 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0812__A2
timestamp 1698175906
transform 1 0 24640 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0812__A3
timestamp 1698175906
transform 1 0 27216 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0815__A2
timestamp 1698175906
transform -1 0 24416 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0816__A1
timestamp 1698175906
transform 1 0 22624 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0818__A1
timestamp 1698175906
transform -1 0 15120 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0818__A2
timestamp 1698175906
transform -1 0 15008 0 1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0819__A1
timestamp 1698175906
transform 1 0 22512 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0819__A2
timestamp 1698175906
transform 1 0 22064 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0820__A1
timestamp 1698175906
transform 1 0 16800 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0820__A2
timestamp 1698175906
transform -1 0 16576 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0821__B
timestamp 1698175906
transform -1 0 17920 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0821__C
timestamp 1698175906
transform -1 0 17472 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0826__A2
timestamp 1698175906
transform 1 0 19152 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0827__A2
timestamp 1698175906
transform 1 0 16352 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0827__B1
timestamp 1698175906
transform -1 0 16352 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0832__A1
timestamp 1698175906
transform 1 0 10528 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0833__C1
timestamp 1698175906
transform 1 0 19600 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0833__C2
timestamp 1698175906
transform 1 0 21392 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0834__I
timestamp 1698175906
transform 1 0 13664 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0835__A1
timestamp 1698175906
transform 1 0 14224 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0836__A1
timestamp 1698175906
transform -1 0 15232 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0837__I
timestamp 1698175906
transform 1 0 17472 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0842__A2
timestamp 1698175906
transform 1 0 29008 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0843__A1
timestamp 1698175906
transform 1 0 29232 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0843__A2
timestamp 1698175906
transform 1 0 28000 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0847__A2
timestamp 1698175906
transform -1 0 21504 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0848__B1
timestamp 1698175906
transform -1 0 25872 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0848__B2
timestamp 1698175906
transform 1 0 25200 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0850__A1
timestamp 1698175906
transform -1 0 11648 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0850__A2
timestamp 1698175906
transform 1 0 11536 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0851__A2
timestamp 1698175906
transform 1 0 22848 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0852__A2
timestamp 1698175906
transform 1 0 12768 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0852__B2
timestamp 1698175906
transform 1 0 12992 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0859__A1
timestamp 1698175906
transform 1 0 20720 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0859__A2
timestamp 1698175906
transform 1 0 21616 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0860__A1
timestamp 1698175906
transform 1 0 27552 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0860__A2
timestamp 1698175906
transform 1 0 23744 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0861__A1
timestamp 1698175906
transform 1 0 27104 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0861__A2
timestamp 1698175906
transform 1 0 26656 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0861__B
timestamp 1698175906
transform -1 0 28784 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0862__A1
timestamp 1698175906
transform 1 0 27216 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0862__B1
timestamp 1698175906
transform 1 0 28784 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0862__B2
timestamp 1698175906
transform 1 0 29232 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0864__A1
timestamp 1698175906
transform 1 0 28672 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0866__B2
timestamp 1698175906
transform 1 0 7280 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0868__A1
timestamp 1698175906
transform -1 0 18144 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0870__A1
timestamp 1698175906
transform 1 0 14560 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0870__A2
timestamp 1698175906
transform 1 0 15008 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0870__B1
timestamp 1698175906
transform 1 0 15456 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0872__I
timestamp 1698175906
transform 1 0 15792 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0875__A1
timestamp 1698175906
transform 1 0 21392 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0876__I
timestamp 1698175906
transform 1 0 26880 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0877__A1
timestamp 1698175906
transform 1 0 18144 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0877__A2
timestamp 1698175906
transform 1 0 19152 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0878__I
timestamp 1698175906
transform -1 0 22288 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0880__A1
timestamp 1698175906
transform 1 0 17472 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0881__I
timestamp 1698175906
transform -1 0 26544 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0883__B1
timestamp 1698175906
transform 1 0 18480 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0883__B2
timestamp 1698175906
transform 1 0 16576 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0893__A2
timestamp 1698175906
transform 1 0 18144 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0894__A1
timestamp 1698175906
transform -1 0 24416 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0894__A2
timestamp 1698175906
transform -1 0 24864 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0896__A1
timestamp 1698175906
transform 1 0 28112 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0897__A2
timestamp 1698175906
transform 1 0 28896 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0898__B1
timestamp 1698175906
transform 1 0 17136 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0899__A2
timestamp 1698175906
transform 1 0 27104 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0899__B
timestamp 1698175906
transform 1 0 27104 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0903__A1
timestamp 1698175906
transform -1 0 7168 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0903__A2
timestamp 1698175906
transform -1 0 6720 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0905__A1
timestamp 1698175906
transform -1 0 12208 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0905__C1
timestamp 1698175906
transform 1 0 13552 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0906__A2
timestamp 1698175906
transform 1 0 12656 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0907__A1
timestamp 1698175906
transform 1 0 15568 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0907__A2
timestamp 1698175906
transform -1 0 14560 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0908__A1
timestamp 1698175906
transform 1 0 14672 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0908__B1
timestamp 1698175906
transform -1 0 15344 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0910__A2
timestamp 1698175906
transform 1 0 22960 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0910__A3
timestamp 1698175906
transform 1 0 22512 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0910__A4
timestamp 1698175906
transform 1 0 22512 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0914__A1
timestamp 1698175906
transform 1 0 24528 0 -1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0919__A1
timestamp 1698175906
transform -1 0 23744 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0919__A2
timestamp 1698175906
transform -1 0 23296 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0920__A1
timestamp 1698175906
transform 1 0 24192 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0921__A2
timestamp 1698175906
transform 1 0 25312 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0922__A1
timestamp 1698175906
transform 1 0 24640 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0923__A1
timestamp 1698175906
transform 1 0 16800 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0924__A1
timestamp 1698175906
transform 1 0 23856 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0924__A2
timestamp 1698175906
transform -1 0 25984 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0928__A1
timestamp 1698175906
transform 1 0 11088 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0928__A2
timestamp 1698175906
transform 1 0 10080 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0929__A1
timestamp 1698175906
transform -1 0 8960 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0930__B1
timestamp 1698175906
transform 1 0 11536 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0930__B2
timestamp 1698175906
transform 1 0 12208 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0931__A1
timestamp 1698175906
transform -1 0 11984 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0932__A2
timestamp 1698175906
transform 1 0 7056 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0934__A2
timestamp 1698175906
transform 1 0 7504 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0937__I
timestamp 1698175906
transform 1 0 14112 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0938__I
timestamp 1698175906
transform 1 0 21840 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0939__A2
timestamp 1698175906
transform 1 0 10528 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0939__B
timestamp 1698175906
transform 1 0 10080 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0940__A1
timestamp 1698175906
transform 1 0 10528 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0940__B
timestamp 1698175906
transform 1 0 10976 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0941__A1
timestamp 1698175906
transform 1 0 4704 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0942__A1
timestamp 1698175906
transform -1 0 4928 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0950__A3
timestamp 1698175906
transform 1 0 23072 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0953__I
timestamp 1698175906
transform 1 0 27440 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0954__A2
timestamp 1698175906
transform -1 0 23184 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0955__A1
timestamp 1698175906
transform 1 0 23184 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0955__A2
timestamp 1698175906
transform 1 0 19824 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0957__A1
timestamp 1698175906
transform 1 0 19264 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0957__B
timestamp 1698175906
transform 1 0 17920 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0959__B2
timestamp 1698175906
transform 1 0 15008 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0960__A1
timestamp 1698175906
transform 1 0 15456 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0961__A1
timestamp 1698175906
transform 1 0 3360 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0961__A3
timestamp 1698175906
transform 1 0 4368 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0967__A1
timestamp 1698175906
transform 1 0 29232 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0974__A1
timestamp 1698175906
transform 1 0 29232 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0974__A2
timestamp 1698175906
transform 1 0 24640 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0976__A2
timestamp 1698175906
transform -1 0 20384 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0977__A1
timestamp 1698175906
transform 1 0 19488 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0979__A2
timestamp 1698175906
transform -1 0 10752 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0980__A1
timestamp 1698175906
transform -1 0 9184 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0980__A2
timestamp 1698175906
transform 1 0 10640 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0980__B1
timestamp 1698175906
transform -1 0 8736 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0981__A1
timestamp 1698175906
transform 1 0 4816 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0981__C2
timestamp 1698175906
transform 1 0 4592 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0983__A4
timestamp 1698175906
transform 1 0 27888 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0986__A1
timestamp 1698175906
transform -1 0 17248 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0987__A1
timestamp 1698175906
transform -1 0 14224 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0988__A3
timestamp 1698175906
transform -1 0 20272 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0989__A1
timestamp 1698175906
transform -1 0 16800 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0989__B
timestamp 1698175906
transform -1 0 18704 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0990__A1
timestamp 1698175906
transform -1 0 15680 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0991__B1
timestamp 1698175906
transform 1 0 13664 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0991__B2
timestamp 1698175906
transform -1 0 16240 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0992__A1
timestamp 1698175906
transform -1 0 15680 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0994__A1
timestamp 1698175906
transform 1 0 22400 0 -1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0995__A3
timestamp 1698175906
transform 1 0 22960 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0998__B
timestamp 1698175906
transform 1 0 26544 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0998__C
timestamp 1698175906
transform 1 0 27664 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1001__A1
timestamp 1698175906
transform -1 0 18704 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1002__A3
timestamp 1698175906
transform 1 0 21840 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1003__A1
timestamp 1698175906
transform 1 0 18928 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1003__A2
timestamp 1698175906
transform -1 0 19600 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1003__B2
timestamp 1698175906
transform 1 0 22400 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1005__A1
timestamp 1698175906
transform -1 0 21168 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1009__A1
timestamp 1698175906
transform 1 0 9184 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1012__A1
timestamp 1698175906
transform -1 0 20720 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1012__A3
timestamp 1698175906
transform -1 0 19824 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1012__A4
timestamp 1698175906
transform -1 0 18704 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1013__C2
timestamp 1698175906
transform 1 0 22736 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1014__A3
timestamp 1698175906
transform 1 0 21504 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1017__A1
timestamp 1698175906
transform 1 0 30352 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1021__A1
timestamp 1698175906
transform -1 0 19712 0 1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1023__A1
timestamp 1698175906
transform 1 0 12880 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1024__A1
timestamp 1698175906
transform 1 0 15344 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1031__A1
timestamp 1698175906
transform 1 0 23632 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1034__I
timestamp 1698175906
transform 1 0 10416 0 1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1037__I
timestamp 1698175906
transform 1 0 12768 0 -1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1038__I
timestamp 1698175906
transform 1 0 12432 0 1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1039__A1
timestamp 1698175906
transform -1 0 12656 0 1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1040__A1
timestamp 1698175906
transform -1 0 12096 0 -1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1042__A1
timestamp 1698175906
transform -1 0 11984 0 1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1043__A1
timestamp 1698175906
transform 1 0 12768 0 1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1045__A1
timestamp 1698175906
transform 1 0 11872 0 1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1046__A1
timestamp 1698175906
transform 1 0 11536 0 1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1048__I
timestamp 1698175906
transform -1 0 31584 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1049__A1
timestamp 1698175906
transform -1 0 13888 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1050__A1
timestamp 1698175906
transform 1 0 12320 0 1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1052__I
timestamp 1698175906
transform -1 0 32704 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1053__I
timestamp 1698175906
transform 1 0 34496 0 1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1054__A1
timestamp 1698175906
transform 1 0 36176 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1055__A1
timestamp 1698175906
transform 1 0 34608 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1057__A1
timestamp 1698175906
transform -1 0 34160 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1058__A1
timestamp 1698175906
transform -1 0 34160 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1060__A1
timestamp 1698175906
transform 1 0 33488 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1061__A1
timestamp 1698175906
transform -1 0 36400 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1063__A2
timestamp 1698175906
transform 1 0 32480 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1064__A1
timestamp 1698175906
transform 1 0 35392 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1065__A2
timestamp 1698175906
transform -1 0 14560 0 1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1066__I
timestamp 1698175906
transform -1 0 21952 0 1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1067__I
timestamp 1698175906
transform 1 0 24080 0 -1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1069__I
timestamp 1698175906
transform 1 0 27440 0 -1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1071__A1
timestamp 1698175906
transform 1 0 23408 0 -1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1073__A1
timestamp 1698175906
transform 1 0 25648 0 1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1075__A1
timestamp 1698175906
transform 1 0 21952 0 1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1077__A1
timestamp 1698175906
transform 1 0 27328 0 1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1078__I
timestamp 1698175906
transform 1 0 37744 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1079__I
timestamp 1698175906
transform -1 0 38976 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1080__I
timestamp 1698175906
transform 1 0 38864 0 1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1082__A1
timestamp 1698175906
transform 1 0 40320 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1084__A1
timestamp 1698175906
transform 1 0 39872 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1086__A1
timestamp 1698175906
transform 1 0 38528 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1088__A1
timestamp 1698175906
transform 1 0 40992 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1089__I
timestamp 1698175906
transform 1 0 29232 0 1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1090__I
timestamp 1698175906
transform 1 0 32592 0 1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1091__I
timestamp 1698175906
transform -1 0 38080 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1093__A1
timestamp 1698175906
transform 1 0 28784 0 -1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1095__A1
timestamp 1698175906
transform 1 0 29232 0 -1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1097__A1
timestamp 1698175906
transform 1 0 32480 0 -1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1098__I
timestamp 1698175906
transform 1 0 37744 0 1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1100__A1
timestamp 1698175906
transform 1 0 32816 0 1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1101__I
timestamp 1698175906
transform 1 0 38192 0 -1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1102__I
timestamp 1698175906
transform 1 0 38416 0 -1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1104__A1
timestamp 1698175906
transform 1 0 38416 0 -1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1106__A1
timestamp 1698175906
transform 1 0 40992 0 -1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1108__A1
timestamp 1698175906
transform 1 0 40992 0 -1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1110__A1
timestamp 1698175906
transform 1 0 40320 0 -1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1114__I
timestamp 1698175906
transform 1 0 16016 0 1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1116__A1
timestamp 1698175906
transform 1 0 15456 0 1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1118__A1
timestamp 1698175906
transform 1 0 15344 0 -1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1120__A1
timestamp 1698175906
transform 1 0 18144 0 1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1122__A1
timestamp 1698175906
transform 1 0 19040 0 -1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1125__I
timestamp 1698175906
transform 1 0 32816 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1127__A1
timestamp 1698175906
transform -1 0 32704 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1129__A1
timestamp 1698175906
transform 1 0 35392 0 -1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1131__A1
timestamp 1698175906
transform 1 0 35728 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1133__A1
timestamp 1698175906
transform 1 0 32144 0 -1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1134__CLK
timestamp 1698175906
transform 1 0 5040 0 -1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1135__CLK
timestamp 1698175906
transform 1 0 5040 0 1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1136__CLK
timestamp 1698175906
transform 1 0 8960 0 1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1137__CLK
timestamp 1698175906
transform 1 0 7616 0 -1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1146__CLK
timestamp 1698175906
transform -1 0 40096 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1150__CLK
timestamp 1698175906
transform 1 0 33152 0 1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1152__CLK
timestamp 1698175906
transform 1 0 37744 0 1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1153__CLK
timestamp 1698175906
transform 1 0 37072 0 1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1154__CLK
timestamp 1698175906
transform 1 0 40432 0 1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1155__CLK
timestamp 1698175906
transform 1 0 41552 0 -1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1156__CLK
timestamp 1698175906
transform 1 0 40880 0 1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1157__CLK
timestamp 1698175906
transform 1 0 39872 0 1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1158__CLK
timestamp 1698175906
transform 1 0 16800 0 1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1159__CLK
timestamp 1698175906
transform 1 0 16464 0 1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1160__CLK
timestamp 1698175906
transform 1 0 21392 0 1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1162__CLK
timestamp 1698175906
transform 1 0 32928 0 1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1163__CLK
timestamp 1698175906
transform 1 0 37072 0 1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1165__CLK
timestamp 1698175906
transform 1 0 32368 0 1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_clkbuf_0_wb_clk_i_I
timestamp 1698175906
transform 1 0 24640 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_clkbuf_2_0__f_wb_clk_i_I
timestamp 1698175906
transform 1 0 27664 0 1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_clkbuf_2_1__f_wb_clk_i_I
timestamp 1698175906
transform 1 0 23072 0 -1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_clkbuf_2_2__f_wb_clk_i_I
timestamp 1698175906
transform 1 0 33712 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_clkbuf_2_3__f_wb_clk_i_I
timestamp 1698175906
transform 1 0 33264 0 -1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input1_I
timestamp 1698175906
transform -1 0 7504 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input2_I
timestamp 1698175906
transform -1 0 23184 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input3_I
timestamp 1698175906
transform -1 0 25424 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input4_I
timestamp 1698175906
transform -1 0 28000 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input5_I
timestamp 1698175906
transform -1 0 29904 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input6_I
timestamp 1698175906
transform -1 0 31808 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input7_I
timestamp 1698175906
transform -1 0 34384 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input8_I
timestamp 1698175906
transform -1 0 36624 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input9_I
timestamp 1698175906
transform -1 0 39424 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input10_I
timestamp 1698175906
transform -1 0 16576 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input11_I
timestamp 1698175906
transform -1 0 18704 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input12_I
timestamp 1698175906
transform -1 0 20384 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input13_I
timestamp 1698175906
transform -1 0 11984 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input14_I
timestamp 1698175906
transform -1 0 9744 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input15_I
timestamp 1698175906
transform 1 0 1792 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input16_I
timestamp 1698175906
transform 1 0 2464 0 1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input17_I
timestamp 1698175906
transform 1 0 2464 0 -1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input18_I
timestamp 1698175906
transform 1 0 2464 0 -1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input19_I
timestamp 1698175906
transform 1 0 2464 0 -1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input20_I
timestamp 1698175906
transform 1 0 3136 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input21_I
timestamp 1698175906
transform -1 0 2240 0 1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input22_I
timestamp 1698175906
transform 1 0 2464 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input23_I
timestamp 1698175906
transform 1 0 1792 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input24_I
timestamp 1698175906
transform 1 0 3136 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input25_I
timestamp 1698175906
transform 1 0 1792 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input26_I
timestamp 1698175906
transform 1 0 2464 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input27_I
timestamp 1698175906
transform 1 0 1792 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input28_I
timestamp 1698175906
transform 1 0 1792 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input29_I
timestamp 1698175906
transform 1 0 2464 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input30_I
timestamp 1698175906
transform 1 0 2464 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input31_I
timestamp 1698175906
transform 1 0 2688 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input32_I
timestamp 1698175906
transform 1 0 2464 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input33_I
timestamp 1698175906
transform 1 0 2464 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input34_I
timestamp 1698175906
transform 1 0 2464 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input35_I
timestamp 1698175906
transform 1 0 2464 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input36_I
timestamp 1698175906
transform 1 0 2464 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input37_I
timestamp 1698175906
transform 1 0 3136 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input38_I
timestamp 1698175906
transform 1 0 2464 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input39_I
timestamp 1698175906
transform 1 0 1792 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input40_I
timestamp 1698175906
transform 1 0 2464 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input41_I
timestamp 1698175906
transform 1 0 2464 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input42_I
timestamp 1698175906
transform 1 0 2464 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input43_I
timestamp 1698175906
transform 1 0 2464 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input44_I
timestamp 1698175906
transform 1 0 2464 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input45_I
timestamp 1698175906
transform 1 0 2464 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input46_I
timestamp 1698175906
transform 1 0 2464 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input47_I
timestamp 1698175906
transform -1 0 14224 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input48_I
timestamp 1698175906
transform -1 0 5152 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output49_I
timestamp 1698175906
transform -1 0 38976 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output50_I
timestamp 1698175906
transform 1 0 43568 0 1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output51_I
timestamp 1698175906
transform 1 0 45360 0 1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output52_I
timestamp 1698175906
transform -1 0 47824 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output53_I
timestamp 1698175906
transform 1 0 50848 0 1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output54_I
timestamp 1698175906
transform 1 0 52080 0 1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output55_I
timestamp 1698175906
transform -1 0 54656 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output56_I
timestamp 1698175906
transform 1 0 55216 0 -1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_16  clkbuf_0_wb_clk_i $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 25088 0 -1 47040
box -86 -86 5686 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_16  clkbuf_2_0__f_wb_clk_i
timestamp 1698175906
transform -1 0 27440 0 1 51744
box -86 -86 5686 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_16  clkbuf_2_1__f_wb_clk_i
timestamp 1698175906
transform -1 0 22848 0 -1 50176
box -86 -86 5686 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_16  clkbuf_2_2__f_wb_clk_i
timestamp 1698175906
transform 1 0 33712 0 -1 45472
box -86 -86 5686 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_16  clkbuf_2_3__f_wb_clk_i
timestamp 1698175906
transform 1 0 33488 0 -1 48608
box -86 -86 5686 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_0_10 $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 2464 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_0_14 $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 2912 0 1 3136
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_0_30 $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 4704 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_0_36 $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 5376 0 1 3136
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_0_70
timestamp 1698175906
transform 1 0 9184 0 1 3136
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_0_104
timestamp 1698175906
transform 1 0 12992 0 1 3136
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_0_138
timestamp 1698175906
transform 1 0 16800 0 1 3136
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_0_172
timestamp 1698175906
transform 1 0 20608 0 1 3136
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_0_206
timestamp 1698175906
transform 1 0 24416 0 1 3136
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_0_240
timestamp 1698175906
transform 1 0 28224 0 1 3136
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_0_274
timestamp 1698175906
transform 1 0 32032 0 1 3136
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_0_308
timestamp 1698175906
transform 1 0 35840 0 1 3136
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_0_342
timestamp 1698175906
transform 1 0 39648 0 1 3136
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_0_376
timestamp 1698175906
transform 1 0 43456 0 1 3136
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_0_410
timestamp 1698175906
transform 1 0 47264 0 1 3136
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_0_444
timestamp 1698175906
transform 1 0 51072 0 1 3136
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_0_478
timestamp 1698175906
transform 1 0 54880 0 1 3136
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_0_494 $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 56672 0 1 3136
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_0_502
timestamp 1698175906
transform 1 0 57568 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_0_506
timestamp 1698175906
transform 1 0 58016 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_0_508 $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 58240 0 1 3136
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_1_8
timestamp 1698175906
transform 1 0 2240 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_1_12
timestamp 1698175906
transform 1 0 2688 0 -1 4704
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_1_44
timestamp 1698175906
transform 1 0 6272 0 -1 4704
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_1_60
timestamp 1698175906
transform 1 0 8064 0 -1 4704
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_1_68
timestamp 1698175906
transform 1 0 8960 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_1_72 $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 9408 0 -1 4704
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_1_136
timestamp 1698175906
transform 1 0 16576 0 -1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_1_142
timestamp 1698175906
transform 1 0 17248 0 -1 4704
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_1_206
timestamp 1698175906
transform 1 0 24416 0 -1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_1_212
timestamp 1698175906
transform 1 0 25088 0 -1 4704
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_1_276
timestamp 1698175906
transform 1 0 32256 0 -1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_1_282
timestamp 1698175906
transform 1 0 32928 0 -1 4704
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_1_346
timestamp 1698175906
transform 1 0 40096 0 -1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_1_352
timestamp 1698175906
transform 1 0 40768 0 -1 4704
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_1_416
timestamp 1698175906
transform 1 0 47936 0 -1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_1_422
timestamp 1698175906
transform 1 0 48608 0 -1 4704
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_1_486
timestamp 1698175906
transform 1 0 55776 0 -1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_1_492
timestamp 1698175906
transform 1 0 56448 0 -1 4704
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_1_508
timestamp 1698175906
transform 1 0 58240 0 -1 4704
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_2_2
timestamp 1698175906
transform 1 0 1568 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_2_6
timestamp 1698175906
transform 1 0 2016 0 1 4704
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_2_22
timestamp 1698175906
transform 1 0 3808 0 1 4704
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_2_30
timestamp 1698175906
transform 1 0 4704 0 1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_2_34
timestamp 1698175906
transform 1 0 5152 0 1 4704
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_2_37
timestamp 1698175906
transform 1 0 5488 0 1 4704
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_2_101
timestamp 1698175906
transform 1 0 12656 0 1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_2_107
timestamp 1698175906
transform 1 0 13328 0 1 4704
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_2_171
timestamp 1698175906
transform 1 0 20496 0 1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_2_177
timestamp 1698175906
transform 1 0 21168 0 1 4704
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_2_241
timestamp 1698175906
transform 1 0 28336 0 1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_2_247
timestamp 1698175906
transform 1 0 29008 0 1 4704
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_2_311
timestamp 1698175906
transform 1 0 36176 0 1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_2_317
timestamp 1698175906
transform 1 0 36848 0 1 4704
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_2_381
timestamp 1698175906
transform 1 0 44016 0 1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_2_387
timestamp 1698175906
transform 1 0 44688 0 1 4704
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_2_451
timestamp 1698175906
transform 1 0 51856 0 1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_2_457
timestamp 1698175906
transform 1 0 52528 0 1 4704
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_2_489
timestamp 1698175906
transform 1 0 56112 0 1 4704
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_2_505
timestamp 1698175906
transform 1 0 57904 0 1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_3_10
timestamp 1698175906
transform 1 0 2464 0 -1 6272
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_3_42
timestamp 1698175906
transform 1 0 6048 0 -1 6272
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_3_58
timestamp 1698175906
transform 1 0 7840 0 -1 6272
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_3_66
timestamp 1698175906
transform 1 0 8736 0 -1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_3_72
timestamp 1698175906
transform 1 0 9408 0 -1 6272
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_3_136
timestamp 1698175906
transform 1 0 16576 0 -1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_3_142
timestamp 1698175906
transform 1 0 17248 0 -1 6272
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_3_206
timestamp 1698175906
transform 1 0 24416 0 -1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_3_212
timestamp 1698175906
transform 1 0 25088 0 -1 6272
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_3_276
timestamp 1698175906
transform 1 0 32256 0 -1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_3_282
timestamp 1698175906
transform 1 0 32928 0 -1 6272
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_3_346
timestamp 1698175906
transform 1 0 40096 0 -1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_3_352
timestamp 1698175906
transform 1 0 40768 0 -1 6272
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_3_416
timestamp 1698175906
transform 1 0 47936 0 -1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_3_422
timestamp 1698175906
transform 1 0 48608 0 -1 6272
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_3_486
timestamp 1698175906
transform 1 0 55776 0 -1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_3_492
timestamp 1698175906
transform 1 0 56448 0 -1 6272
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_3_508
timestamp 1698175906
transform 1 0 58240 0 -1 6272
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_4_2
timestamp 1698175906
transform 1 0 1568 0 1 6272
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_4_34
timestamp 1698175906
transform 1 0 5152 0 1 6272
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_4_37
timestamp 1698175906
transform 1 0 5488 0 1 6272
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_4_101
timestamp 1698175906
transform 1 0 12656 0 1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_4_107
timestamp 1698175906
transform 1 0 13328 0 1 6272
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_4_171
timestamp 1698175906
transform 1 0 20496 0 1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_4_177
timestamp 1698175906
transform 1 0 21168 0 1 6272
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_4_241
timestamp 1698175906
transform 1 0 28336 0 1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_4_247
timestamp 1698175906
transform 1 0 29008 0 1 6272
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_4_311
timestamp 1698175906
transform 1 0 36176 0 1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_4_317
timestamp 1698175906
transform 1 0 36848 0 1 6272
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_4_381
timestamp 1698175906
transform 1 0 44016 0 1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_4_387
timestamp 1698175906
transform 1 0 44688 0 1 6272
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_4_451
timestamp 1698175906
transform 1 0 51856 0 1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_4_457
timestamp 1698175906
transform 1 0 52528 0 1 6272
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_4_489
timestamp 1698175906
transform 1 0 56112 0 1 6272
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_4_505
timestamp 1698175906
transform 1 0 57904 0 1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_5_2
timestamp 1698175906
transform 1 0 1568 0 -1 7840
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_5_66
timestamp 1698175906
transform 1 0 8736 0 -1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_5_72
timestamp 1698175906
transform 1 0 9408 0 -1 7840
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_5_136
timestamp 1698175906
transform 1 0 16576 0 -1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_5_142
timestamp 1698175906
transform 1 0 17248 0 -1 7840
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_5_206
timestamp 1698175906
transform 1 0 24416 0 -1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_5_212
timestamp 1698175906
transform 1 0 25088 0 -1 7840
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_5_276
timestamp 1698175906
transform 1 0 32256 0 -1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_5_282
timestamp 1698175906
transform 1 0 32928 0 -1 7840
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_5_346
timestamp 1698175906
transform 1 0 40096 0 -1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_5_352
timestamp 1698175906
transform 1 0 40768 0 -1 7840
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_5_416
timestamp 1698175906
transform 1 0 47936 0 -1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_5_422
timestamp 1698175906
transform 1 0 48608 0 -1 7840
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_5_486
timestamp 1698175906
transform 1 0 55776 0 -1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_5_492
timestamp 1698175906
transform 1 0 56448 0 -1 7840
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_5_508
timestamp 1698175906
transform 1 0 58240 0 -1 7840
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_6_8
timestamp 1698175906
transform 1 0 2240 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_6_12
timestamp 1698175906
transform 1 0 2688 0 1 7840
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_6_28
timestamp 1698175906
transform 1 0 4480 0 1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_6_32
timestamp 1698175906
transform 1 0 4928 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_6_34
timestamp 1698175906
transform 1 0 5152 0 1 7840
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_6_37
timestamp 1698175906
transform 1 0 5488 0 1 7840
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_6_101
timestamp 1698175906
transform 1 0 12656 0 1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_6_107
timestamp 1698175906
transform 1 0 13328 0 1 7840
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_6_171
timestamp 1698175906
transform 1 0 20496 0 1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_6_177
timestamp 1698175906
transform 1 0 21168 0 1 7840
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_6_241
timestamp 1698175906
transform 1 0 28336 0 1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_6_247
timestamp 1698175906
transform 1 0 29008 0 1 7840
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_6_311
timestamp 1698175906
transform 1 0 36176 0 1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_6_317
timestamp 1698175906
transform 1 0 36848 0 1 7840
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_6_381
timestamp 1698175906
transform 1 0 44016 0 1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_6_387
timestamp 1698175906
transform 1 0 44688 0 1 7840
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_6_451
timestamp 1698175906
transform 1 0 51856 0 1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_6_457
timestamp 1698175906
transform 1 0 52528 0 1 7840
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_6_489
timestamp 1698175906
transform 1 0 56112 0 1 7840
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_6_505
timestamp 1698175906
transform 1 0 57904 0 1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_7_2
timestamp 1698175906
transform 1 0 1568 0 -1 9408
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_7_66
timestamp 1698175906
transform 1 0 8736 0 -1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_7_72
timestamp 1698175906
transform 1 0 9408 0 -1 9408
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_7_136
timestamp 1698175906
transform 1 0 16576 0 -1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_7_142
timestamp 1698175906
transform 1 0 17248 0 -1 9408
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_7_206
timestamp 1698175906
transform 1 0 24416 0 -1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_7_212
timestamp 1698175906
transform 1 0 25088 0 -1 9408
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_7_276
timestamp 1698175906
transform 1 0 32256 0 -1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_7_282
timestamp 1698175906
transform 1 0 32928 0 -1 9408
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_7_346
timestamp 1698175906
transform 1 0 40096 0 -1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_7_352
timestamp 1698175906
transform 1 0 40768 0 -1 9408
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_7_416
timestamp 1698175906
transform 1 0 47936 0 -1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_7_422
timestamp 1698175906
transform 1 0 48608 0 -1 9408
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_7_486
timestamp 1698175906
transform 1 0 55776 0 -1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_7_492
timestamp 1698175906
transform 1 0 56448 0 -1 9408
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_7_508
timestamp 1698175906
transform 1 0 58240 0 -1 9408
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_8_8
timestamp 1698175906
transform 1 0 2240 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_8_12
timestamp 1698175906
transform 1 0 2688 0 1 9408
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_8_28
timestamp 1698175906
transform 1 0 4480 0 1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_8_32
timestamp 1698175906
transform 1 0 4928 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_8_34
timestamp 1698175906
transform 1 0 5152 0 1 9408
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_8_37
timestamp 1698175906
transform 1 0 5488 0 1 9408
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_8_101
timestamp 1698175906
transform 1 0 12656 0 1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_8_107
timestamp 1698175906
transform 1 0 13328 0 1 9408
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_8_171
timestamp 1698175906
transform 1 0 20496 0 1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_8_177
timestamp 1698175906
transform 1 0 21168 0 1 9408
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_8_241
timestamp 1698175906
transform 1 0 28336 0 1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_8_247
timestamp 1698175906
transform 1 0 29008 0 1 9408
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_8_311
timestamp 1698175906
transform 1 0 36176 0 1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_8_317
timestamp 1698175906
transform 1 0 36848 0 1 9408
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_8_381
timestamp 1698175906
transform 1 0 44016 0 1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_8_387
timestamp 1698175906
transform 1 0 44688 0 1 9408
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_8_451
timestamp 1698175906
transform 1 0 51856 0 1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_8_457
timestamp 1698175906
transform 1 0 52528 0 1 9408
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_8_489
timestamp 1698175906
transform 1 0 56112 0 1 9408
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_8_505
timestamp 1698175906
transform 1 0 57904 0 1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_9_2
timestamp 1698175906
transform 1 0 1568 0 -1 10976
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_9_66
timestamp 1698175906
transform 1 0 8736 0 -1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_9_72
timestamp 1698175906
transform 1 0 9408 0 -1 10976
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_9_136
timestamp 1698175906
transform 1 0 16576 0 -1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_9_142
timestamp 1698175906
transform 1 0 17248 0 -1 10976
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_9_206
timestamp 1698175906
transform 1 0 24416 0 -1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_9_212
timestamp 1698175906
transform 1 0 25088 0 -1 10976
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_9_276
timestamp 1698175906
transform 1 0 32256 0 -1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_9_282
timestamp 1698175906
transform 1 0 32928 0 -1 10976
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_9_346
timestamp 1698175906
transform 1 0 40096 0 -1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_9_352
timestamp 1698175906
transform 1 0 40768 0 -1 10976
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_9_416
timestamp 1698175906
transform 1 0 47936 0 -1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_9_422
timestamp 1698175906
transform 1 0 48608 0 -1 10976
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_9_486
timestamp 1698175906
transform 1 0 55776 0 -1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_9_492
timestamp 1698175906
transform 1 0 56448 0 -1 10976
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_9_508
timestamp 1698175906
transform 1 0 58240 0 -1 10976
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_10_8
timestamp 1698175906
transform 1 0 2240 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_10_12
timestamp 1698175906
transform 1 0 2688 0 1 10976
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_10_28
timestamp 1698175906
transform 1 0 4480 0 1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_10_32
timestamp 1698175906
transform 1 0 4928 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_10_34
timestamp 1698175906
transform 1 0 5152 0 1 10976
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_10_37
timestamp 1698175906
transform 1 0 5488 0 1 10976
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_10_101
timestamp 1698175906
transform 1 0 12656 0 1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_10_107
timestamp 1698175906
transform 1 0 13328 0 1 10976
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_10_171
timestamp 1698175906
transform 1 0 20496 0 1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_10_177
timestamp 1698175906
transform 1 0 21168 0 1 10976
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_10_241
timestamp 1698175906
transform 1 0 28336 0 1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_10_247
timestamp 1698175906
transform 1 0 29008 0 1 10976
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_10_311
timestamp 1698175906
transform 1 0 36176 0 1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_10_317
timestamp 1698175906
transform 1 0 36848 0 1 10976
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_10_381
timestamp 1698175906
transform 1 0 44016 0 1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_10_387
timestamp 1698175906
transform 1 0 44688 0 1 10976
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_10_451
timestamp 1698175906
transform 1 0 51856 0 1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_10_457
timestamp 1698175906
transform 1 0 52528 0 1 10976
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_10_489
timestamp 1698175906
transform 1 0 56112 0 1 10976
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_10_505
timestamp 1698175906
transform 1 0 57904 0 1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_11_2
timestamp 1698175906
transform 1 0 1568 0 -1 12544
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_11_66
timestamp 1698175906
transform 1 0 8736 0 -1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_11_72
timestamp 1698175906
transform 1 0 9408 0 -1 12544
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_11_136
timestamp 1698175906
transform 1 0 16576 0 -1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_11_142
timestamp 1698175906
transform 1 0 17248 0 -1 12544
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_11_206
timestamp 1698175906
transform 1 0 24416 0 -1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_11_212
timestamp 1698175906
transform 1 0 25088 0 -1 12544
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_11_276
timestamp 1698175906
transform 1 0 32256 0 -1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_11_282
timestamp 1698175906
transform 1 0 32928 0 -1 12544
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_11_346
timestamp 1698175906
transform 1 0 40096 0 -1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_11_352
timestamp 1698175906
transform 1 0 40768 0 -1 12544
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_11_416
timestamp 1698175906
transform 1 0 47936 0 -1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_11_422
timestamp 1698175906
transform 1 0 48608 0 -1 12544
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_11_486
timestamp 1698175906
transform 1 0 55776 0 -1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_11_492
timestamp 1698175906
transform 1 0 56448 0 -1 12544
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_11_508
timestamp 1698175906
transform 1 0 58240 0 -1 12544
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_12_8
timestamp 1698175906
transform 1 0 2240 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_12_12
timestamp 1698175906
transform 1 0 2688 0 1 12544
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_12_28
timestamp 1698175906
transform 1 0 4480 0 1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_12_32
timestamp 1698175906
transform 1 0 4928 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_12_34
timestamp 1698175906
transform 1 0 5152 0 1 12544
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_12_37
timestamp 1698175906
transform 1 0 5488 0 1 12544
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_12_101
timestamp 1698175906
transform 1 0 12656 0 1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_12_107
timestamp 1698175906
transform 1 0 13328 0 1 12544
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_12_171
timestamp 1698175906
transform 1 0 20496 0 1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_12_177
timestamp 1698175906
transform 1 0 21168 0 1 12544
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_12_241
timestamp 1698175906
transform 1 0 28336 0 1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_12_247
timestamp 1698175906
transform 1 0 29008 0 1 12544
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_12_311
timestamp 1698175906
transform 1 0 36176 0 1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_12_317
timestamp 1698175906
transform 1 0 36848 0 1 12544
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_12_381
timestamp 1698175906
transform 1 0 44016 0 1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_12_387
timestamp 1698175906
transform 1 0 44688 0 1 12544
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_12_451
timestamp 1698175906
transform 1 0 51856 0 1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_12_457
timestamp 1698175906
transform 1 0 52528 0 1 12544
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_12_489
timestamp 1698175906
transform 1 0 56112 0 1 12544
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_12_505
timestamp 1698175906
transform 1 0 57904 0 1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_13_2
timestamp 1698175906
transform 1 0 1568 0 -1 14112
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_13_66
timestamp 1698175906
transform 1 0 8736 0 -1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_13_72
timestamp 1698175906
transform 1 0 9408 0 -1 14112
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_13_136
timestamp 1698175906
transform 1 0 16576 0 -1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_13_142
timestamp 1698175906
transform 1 0 17248 0 -1 14112
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_13_206
timestamp 1698175906
transform 1 0 24416 0 -1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_13_212
timestamp 1698175906
transform 1 0 25088 0 -1 14112
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_13_276
timestamp 1698175906
transform 1 0 32256 0 -1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_13_282
timestamp 1698175906
transform 1 0 32928 0 -1 14112
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_13_346
timestamp 1698175906
transform 1 0 40096 0 -1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_13_352
timestamp 1698175906
transform 1 0 40768 0 -1 14112
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_13_416
timestamp 1698175906
transform 1 0 47936 0 -1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_13_422
timestamp 1698175906
transform 1 0 48608 0 -1 14112
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_13_486
timestamp 1698175906
transform 1 0 55776 0 -1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_13_492
timestamp 1698175906
transform 1 0 56448 0 -1 14112
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_13_508
timestamp 1698175906
transform 1 0 58240 0 -1 14112
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_14_2
timestamp 1698175906
transform 1 0 1568 0 1 14112
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_14_34
timestamp 1698175906
transform 1 0 5152 0 1 14112
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_14_37
timestamp 1698175906
transform 1 0 5488 0 1 14112
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_14_101
timestamp 1698175906
transform 1 0 12656 0 1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_14_107
timestamp 1698175906
transform 1 0 13328 0 1 14112
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_14_171
timestamp 1698175906
transform 1 0 20496 0 1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_14_177
timestamp 1698175906
transform 1 0 21168 0 1 14112
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_14_241
timestamp 1698175906
transform 1 0 28336 0 1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_14_247
timestamp 1698175906
transform 1 0 29008 0 1 14112
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_14_311
timestamp 1698175906
transform 1 0 36176 0 1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_14_317
timestamp 1698175906
transform 1 0 36848 0 1 14112
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_14_381
timestamp 1698175906
transform 1 0 44016 0 1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_14_387
timestamp 1698175906
transform 1 0 44688 0 1 14112
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_14_451
timestamp 1698175906
transform 1 0 51856 0 1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_14_457
timestamp 1698175906
transform 1 0 52528 0 1 14112
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_14_489
timestamp 1698175906
transform 1 0 56112 0 1 14112
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_14_505
timestamp 1698175906
transform 1 0 57904 0 1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_15_8
timestamp 1698175906
transform 1 0 2240 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_15_12
timestamp 1698175906
transform 1 0 2688 0 -1 15680
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_15_44
timestamp 1698175906
transform 1 0 6272 0 -1 15680
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_15_60
timestamp 1698175906
transform 1 0 8064 0 -1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_15_68
timestamp 1698175906
transform 1 0 8960 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_15_72
timestamp 1698175906
transform 1 0 9408 0 -1 15680
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_15_136
timestamp 1698175906
transform 1 0 16576 0 -1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_15_142
timestamp 1698175906
transform 1 0 17248 0 -1 15680
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_15_206
timestamp 1698175906
transform 1 0 24416 0 -1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_15_212
timestamp 1698175906
transform 1 0 25088 0 -1 15680
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_15_276
timestamp 1698175906
transform 1 0 32256 0 -1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_15_282
timestamp 1698175906
transform 1 0 32928 0 -1 15680
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_15_346
timestamp 1698175906
transform 1 0 40096 0 -1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_15_352
timestamp 1698175906
transform 1 0 40768 0 -1 15680
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_15_416
timestamp 1698175906
transform 1 0 47936 0 -1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_15_422
timestamp 1698175906
transform 1 0 48608 0 -1 15680
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_15_486
timestamp 1698175906
transform 1 0 55776 0 -1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_15_492
timestamp 1698175906
transform 1 0 56448 0 -1 15680
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_15_508
timestamp 1698175906
transform 1 0 58240 0 -1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_16_2
timestamp 1698175906
transform 1 0 1568 0 1 15680
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_16_34
timestamp 1698175906
transform 1 0 5152 0 1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_16_37
timestamp 1698175906
transform 1 0 5488 0 1 15680
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_16_101
timestamp 1698175906
transform 1 0 12656 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_16_107
timestamp 1698175906
transform 1 0 13328 0 1 15680
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_16_171
timestamp 1698175906
transform 1 0 20496 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_16_177
timestamp 1698175906
transform 1 0 21168 0 1 15680
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_16_241
timestamp 1698175906
transform 1 0 28336 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_16_247
timestamp 1698175906
transform 1 0 29008 0 1 15680
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_16_311
timestamp 1698175906
transform 1 0 36176 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_16_317
timestamp 1698175906
transform 1 0 36848 0 1 15680
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_16_381
timestamp 1698175906
transform 1 0 44016 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_16_387
timestamp 1698175906
transform 1 0 44688 0 1 15680
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_16_451
timestamp 1698175906
transform 1 0 51856 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_16_457
timestamp 1698175906
transform 1 0 52528 0 1 15680
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_16_489
timestamp 1698175906
transform 1 0 56112 0 1 15680
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_16_505
timestamp 1698175906
transform 1 0 57904 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_17_8
timestamp 1698175906
transform 1 0 2240 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_17_12
timestamp 1698175906
transform 1 0 2688 0 -1 17248
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_17_44
timestamp 1698175906
transform 1 0 6272 0 -1 17248
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_17_60
timestamp 1698175906
transform 1 0 8064 0 -1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_17_68
timestamp 1698175906
transform 1 0 8960 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_17_72
timestamp 1698175906
transform 1 0 9408 0 -1 17248
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_17_136
timestamp 1698175906
transform 1 0 16576 0 -1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_17_142
timestamp 1698175906
transform 1 0 17248 0 -1 17248
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_17_206
timestamp 1698175906
transform 1 0 24416 0 -1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_17_212
timestamp 1698175906
transform 1 0 25088 0 -1 17248
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_17_276
timestamp 1698175906
transform 1 0 32256 0 -1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_17_282
timestamp 1698175906
transform 1 0 32928 0 -1 17248
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_17_346
timestamp 1698175906
transform 1 0 40096 0 -1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_17_352
timestamp 1698175906
transform 1 0 40768 0 -1 17248
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_17_416
timestamp 1698175906
transform 1 0 47936 0 -1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_17_422
timestamp 1698175906
transform 1 0 48608 0 -1 17248
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_17_486
timestamp 1698175906
transform 1 0 55776 0 -1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_17_492
timestamp 1698175906
transform 1 0 56448 0 -1 17248
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_17_508
timestamp 1698175906
transform 1 0 58240 0 -1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_18_2
timestamp 1698175906
transform 1 0 1568 0 1 17248
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_18_34
timestamp 1698175906
transform 1 0 5152 0 1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_18_37
timestamp 1698175906
transform 1 0 5488 0 1 17248
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_18_101
timestamp 1698175906
transform 1 0 12656 0 1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_18_107
timestamp 1698175906
transform 1 0 13328 0 1 17248
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_18_171
timestamp 1698175906
transform 1 0 20496 0 1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_18_177
timestamp 1698175906
transform 1 0 21168 0 1 17248
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_18_241
timestamp 1698175906
transform 1 0 28336 0 1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_18_247
timestamp 1698175906
transform 1 0 29008 0 1 17248
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_18_311
timestamp 1698175906
transform 1 0 36176 0 1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_18_317
timestamp 1698175906
transform 1 0 36848 0 1 17248
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_18_381
timestamp 1698175906
transform 1 0 44016 0 1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_18_387
timestamp 1698175906
transform 1 0 44688 0 1 17248
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_18_451
timestamp 1698175906
transform 1 0 51856 0 1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_18_457
timestamp 1698175906
transform 1 0 52528 0 1 17248
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_18_489
timestamp 1698175906
transform 1 0 56112 0 1 17248
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_18_505
timestamp 1698175906
transform 1 0 57904 0 1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_19_8
timestamp 1698175906
transform 1 0 2240 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_19_12
timestamp 1698175906
transform 1 0 2688 0 -1 18816
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_19_44
timestamp 1698175906
transform 1 0 6272 0 -1 18816
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_19_60
timestamp 1698175906
transform 1 0 8064 0 -1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_19_68
timestamp 1698175906
transform 1 0 8960 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_19_72
timestamp 1698175906
transform 1 0 9408 0 -1 18816
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_19_136
timestamp 1698175906
transform 1 0 16576 0 -1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_19_142
timestamp 1698175906
transform 1 0 17248 0 -1 18816
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_19_206
timestamp 1698175906
transform 1 0 24416 0 -1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_19_212
timestamp 1698175906
transform 1 0 25088 0 -1 18816
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_19_276
timestamp 1698175906
transform 1 0 32256 0 -1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_19_282
timestamp 1698175906
transform 1 0 32928 0 -1 18816
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_19_346
timestamp 1698175906
transform 1 0 40096 0 -1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_19_352
timestamp 1698175906
transform 1 0 40768 0 -1 18816
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_19_416
timestamp 1698175906
transform 1 0 47936 0 -1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_19_422
timestamp 1698175906
transform 1 0 48608 0 -1 18816
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_19_486
timestamp 1698175906
transform 1 0 55776 0 -1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_19_492
timestamp 1698175906
transform 1 0 56448 0 -1 18816
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_19_508
timestamp 1698175906
transform 1 0 58240 0 -1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_20_2
timestamp 1698175906
transform 1 0 1568 0 1 18816
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_20_34
timestamp 1698175906
transform 1 0 5152 0 1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_20_37
timestamp 1698175906
transform 1 0 5488 0 1 18816
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_20_101
timestamp 1698175906
transform 1 0 12656 0 1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_20_107
timestamp 1698175906
transform 1 0 13328 0 1 18816
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_20_171
timestamp 1698175906
transform 1 0 20496 0 1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_20_177
timestamp 1698175906
transform 1 0 21168 0 1 18816
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_20_241
timestamp 1698175906
transform 1 0 28336 0 1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_20_247
timestamp 1698175906
transform 1 0 29008 0 1 18816
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_20_311
timestamp 1698175906
transform 1 0 36176 0 1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_20_317
timestamp 1698175906
transform 1 0 36848 0 1 18816
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_20_381
timestamp 1698175906
transform 1 0 44016 0 1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_20_387
timestamp 1698175906
transform 1 0 44688 0 1 18816
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_20_451
timestamp 1698175906
transform 1 0 51856 0 1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_20_457
timestamp 1698175906
transform 1 0 52528 0 1 18816
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_20_489
timestamp 1698175906
transform 1 0 56112 0 1 18816
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_20_505
timestamp 1698175906
transform 1 0 57904 0 1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_21_2
timestamp 1698175906
transform 1 0 1568 0 -1 20384
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_21_66
timestamp 1698175906
transform 1 0 8736 0 -1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_21_72
timestamp 1698175906
transform 1 0 9408 0 -1 20384
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_21_136
timestamp 1698175906
transform 1 0 16576 0 -1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_21_142
timestamp 1698175906
transform 1 0 17248 0 -1 20384
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_21_206
timestamp 1698175906
transform 1 0 24416 0 -1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_21_212
timestamp 1698175906
transform 1 0 25088 0 -1 20384
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_21_276
timestamp 1698175906
transform 1 0 32256 0 -1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_21_282
timestamp 1698175906
transform 1 0 32928 0 -1 20384
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_21_346
timestamp 1698175906
transform 1 0 40096 0 -1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_21_352
timestamp 1698175906
transform 1 0 40768 0 -1 20384
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_21_416
timestamp 1698175906
transform 1 0 47936 0 -1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_21_422
timestamp 1698175906
transform 1 0 48608 0 -1 20384
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_21_486
timestamp 1698175906
transform 1 0 55776 0 -1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_21_492
timestamp 1698175906
transform 1 0 56448 0 -1 20384
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_21_508
timestamp 1698175906
transform 1 0 58240 0 -1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_22_8
timestamp 1698175906
transform 1 0 2240 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_22_12
timestamp 1698175906
transform 1 0 2688 0 1 20384
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_22_28
timestamp 1698175906
transform 1 0 4480 0 1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_22_32
timestamp 1698175906
transform 1 0 4928 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_22_34
timestamp 1698175906
transform 1 0 5152 0 1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_22_37
timestamp 1698175906
transform 1 0 5488 0 1 20384
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_22_101
timestamp 1698175906
transform 1 0 12656 0 1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_22_107
timestamp 1698175906
transform 1 0 13328 0 1 20384
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_22_171
timestamp 1698175906
transform 1 0 20496 0 1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_22_177
timestamp 1698175906
transform 1 0 21168 0 1 20384
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_22_241
timestamp 1698175906
transform 1 0 28336 0 1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_22_247
timestamp 1698175906
transform 1 0 29008 0 1 20384
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_22_311
timestamp 1698175906
transform 1 0 36176 0 1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_22_317
timestamp 1698175906
transform 1 0 36848 0 1 20384
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_22_381
timestamp 1698175906
transform 1 0 44016 0 1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_22_387
timestamp 1698175906
transform 1 0 44688 0 1 20384
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_22_451
timestamp 1698175906
transform 1 0 51856 0 1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_22_457
timestamp 1698175906
transform 1 0 52528 0 1 20384
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_22_489
timestamp 1698175906
transform 1 0 56112 0 1 20384
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_22_505
timestamp 1698175906
transform 1 0 57904 0 1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_23_2
timestamp 1698175906
transform 1 0 1568 0 -1 21952
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_23_66
timestamp 1698175906
transform 1 0 8736 0 -1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_23_72
timestamp 1698175906
transform 1 0 9408 0 -1 21952
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_23_136
timestamp 1698175906
transform 1 0 16576 0 -1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_23_142
timestamp 1698175906
transform 1 0 17248 0 -1 21952
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_23_206
timestamp 1698175906
transform 1 0 24416 0 -1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_23_212
timestamp 1698175906
transform 1 0 25088 0 -1 21952
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_23_276
timestamp 1698175906
transform 1 0 32256 0 -1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_23_282
timestamp 1698175906
transform 1 0 32928 0 -1 21952
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_23_346
timestamp 1698175906
transform 1 0 40096 0 -1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_23_352
timestamp 1698175906
transform 1 0 40768 0 -1 21952
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_23_416
timestamp 1698175906
transform 1 0 47936 0 -1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_23_422
timestamp 1698175906
transform 1 0 48608 0 -1 21952
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_23_486
timestamp 1698175906
transform 1 0 55776 0 -1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_23_492
timestamp 1698175906
transform 1 0 56448 0 -1 21952
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_23_508
timestamp 1698175906
transform 1 0 58240 0 -1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_24_8
timestamp 1698175906
transform 1 0 2240 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_24_12
timestamp 1698175906
transform 1 0 2688 0 1 21952
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_24_28
timestamp 1698175906
transform 1 0 4480 0 1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_24_32
timestamp 1698175906
transform 1 0 4928 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_24_34
timestamp 1698175906
transform 1 0 5152 0 1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_24_37
timestamp 1698175906
transform 1 0 5488 0 1 21952
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_24_101
timestamp 1698175906
transform 1 0 12656 0 1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_24_107
timestamp 1698175906
transform 1 0 13328 0 1 21952
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_24_123
timestamp 1698175906
transform 1 0 15120 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_24_125
timestamp 1698175906
transform 1 0 15344 0 1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_24_128
timestamp 1698175906
transform 1 0 15680 0 1 21952
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_24_160
timestamp 1698175906
transform 1 0 19264 0 1 21952
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_24_168
timestamp 1698175906
transform 1 0 20160 0 1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_24_172
timestamp 1698175906
transform 1 0 20608 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_24_174
timestamp 1698175906
transform 1 0 20832 0 1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_24_177
timestamp 1698175906
transform 1 0 21168 0 1 21952
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_24_241
timestamp 1698175906
transform 1 0 28336 0 1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_24_247
timestamp 1698175906
transform 1 0 29008 0 1 21952
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_24_311
timestamp 1698175906
transform 1 0 36176 0 1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_24_317
timestamp 1698175906
transform 1 0 36848 0 1 21952
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_24_381
timestamp 1698175906
transform 1 0 44016 0 1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_24_387
timestamp 1698175906
transform 1 0 44688 0 1 21952
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_24_451
timestamp 1698175906
transform 1 0 51856 0 1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_24_457
timestamp 1698175906
transform 1 0 52528 0 1 21952
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_24_489
timestamp 1698175906
transform 1 0 56112 0 1 21952
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_24_505
timestamp 1698175906
transform 1 0 57904 0 1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_25_2
timestamp 1698175906
transform 1 0 1568 0 -1 23520
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_25_66
timestamp 1698175906
transform 1 0 8736 0 -1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_25_72
timestamp 1698175906
transform 1 0 9408 0 -1 23520
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_25_104
timestamp 1698175906
transform 1 0 12992 0 -1 23520
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_25_120
timestamp 1698175906
transform 1 0 14784 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_25_124
timestamp 1698175906
transform 1 0 15232 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_25_133
timestamp 1698175906
transform 1 0 16240 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_25_135
timestamp 1698175906
transform 1 0 16464 0 -1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_25_138
timestamp 1698175906
transform 1 0 16800 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_25_142
timestamp 1698175906
transform 1 0 17248 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_25_146
timestamp 1698175906
transform 1 0 17696 0 -1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_25_150
timestamp 1698175906
transform 1 0 18144 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_25_152
timestamp 1698175906
transform 1 0 18368 0 -1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_25_155
timestamp 1698175906
transform 1 0 18704 0 -1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_25_161
timestamp 1698175906
transform 1 0 19376 0 -1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_25_169
timestamp 1698175906
transform 1 0 20272 0 -1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_25_173
timestamp 1698175906
transform 1 0 20720 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_25_183
timestamp 1698175906
transform 1 0 21840 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_25_187
timestamp 1698175906
transform 1 0 22288 0 -1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_25_191
timestamp 1698175906
transform 1 0 22736 0 -1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_25_194
timestamp 1698175906
transform 1 0 23072 0 -1 23520
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_25_212
timestamp 1698175906
transform 1 0 25088 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_25_216
timestamp 1698175906
transform 1 0 25536 0 -1 23520
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_25_282
timestamp 1698175906
transform 1 0 32928 0 -1 23520
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_25_346
timestamp 1698175906
transform 1 0 40096 0 -1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_25_352
timestamp 1698175906
transform 1 0 40768 0 -1 23520
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_25_416
timestamp 1698175906
transform 1 0 47936 0 -1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_25_422
timestamp 1698175906
transform 1 0 48608 0 -1 23520
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_25_486
timestamp 1698175906
transform 1 0 55776 0 -1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_25_492
timestamp 1698175906
transform 1 0 56448 0 -1 23520
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_25_508
timestamp 1698175906
transform 1 0 58240 0 -1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_26_8
timestamp 1698175906
transform 1 0 2240 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_26_12
timestamp 1698175906
transform 1 0 2688 0 1 23520
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_26_28
timestamp 1698175906
transform 1 0 4480 0 1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_26_32
timestamp 1698175906
transform 1 0 4928 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_26_34
timestamp 1698175906
transform 1 0 5152 0 1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_26_37
timestamp 1698175906
transform 1 0 5488 0 1 23520
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_26_69
timestamp 1698175906
transform 1 0 9072 0 1 23520
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_26_85
timestamp 1698175906
transform 1 0 10864 0 1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_26_89
timestamp 1698175906
transform 1 0 11312 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_26_93
timestamp 1698175906
transform 1 0 11760 0 1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_26_101
timestamp 1698175906
transform 1 0 12656 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_26_129
timestamp 1698175906
transform 1 0 15792 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_26_192
timestamp 1698175906
transform 1 0 22848 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_26_194
timestamp 1698175906
transform 1 0 23072 0 1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_26_211
timestamp 1698175906
transform 1 0 24976 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_26_215
timestamp 1698175906
transform 1 0 25424 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_26_219
timestamp 1698175906
transform 1 0 25872 0 1 23520
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_26_235
timestamp 1698175906
transform 1 0 27664 0 1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_26_243
timestamp 1698175906
transform 1 0 28560 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_26_247
timestamp 1698175906
transform 1 0 29008 0 1 23520
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_26_311
timestamp 1698175906
transform 1 0 36176 0 1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_26_317
timestamp 1698175906
transform 1 0 36848 0 1 23520
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_26_381
timestamp 1698175906
transform 1 0 44016 0 1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_26_387
timestamp 1698175906
transform 1 0 44688 0 1 23520
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_26_451
timestamp 1698175906
transform 1 0 51856 0 1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_26_457
timestamp 1698175906
transform 1 0 52528 0 1 23520
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_26_489
timestamp 1698175906
transform 1 0 56112 0 1 23520
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_26_505
timestamp 1698175906
transform 1 0 57904 0 1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_27_2
timestamp 1698175906
transform 1 0 1568 0 -1 25088
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_27_34
timestamp 1698175906
transform 1 0 5152 0 -1 25088
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_27_42
timestamp 1698175906
transform 1 0 6048 0 -1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_27_46
timestamp 1698175906
transform 1 0 6496 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_27_48
timestamp 1698175906
transform 1 0 6720 0 -1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_27_59
timestamp 1698175906
transform 1 0 7952 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_27_63
timestamp 1698175906
transform 1 0 8400 0 -1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_27_67
timestamp 1698175906
transform 1 0 8848 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_27_69
timestamp 1698175906
transform 1 0 9072 0 -1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_27_72
timestamp 1698175906
transform 1 0 9408 0 -1 25088
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_27_80
timestamp 1698175906
transform 1 0 10304 0 -1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_27_84
timestamp 1698175906
transform 1 0 10752 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_27_86
timestamp 1698175906
transform 1 0 10976 0 -1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_27_89
timestamp 1698175906
transform 1 0 11312 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_27_142
timestamp 1698175906
transform 1 0 17248 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_27_220
timestamp 1698175906
transform 1 0 25984 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_27_224
timestamp 1698175906
transform 1 0 26432 0 -1 25088
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_27_256
timestamp 1698175906
transform 1 0 30016 0 -1 25088
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_27_272
timestamp 1698175906
transform 1 0 31808 0 -1 25088
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_27_282
timestamp 1698175906
transform 1 0 32928 0 -1 25088
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_27_346
timestamp 1698175906
transform 1 0 40096 0 -1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_27_352
timestamp 1698175906
transform 1 0 40768 0 -1 25088
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_27_416
timestamp 1698175906
transform 1 0 47936 0 -1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_27_422
timestamp 1698175906
transform 1 0 48608 0 -1 25088
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_27_486
timestamp 1698175906
transform 1 0 55776 0 -1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_27_492
timestamp 1698175906
transform 1 0 56448 0 -1 25088
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_27_508
timestamp 1698175906
transform 1 0 58240 0 -1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_28_8
timestamp 1698175906
transform 1 0 2240 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_28_12
timestamp 1698175906
transform 1 0 2688 0 1 25088
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_28_28
timestamp 1698175906
transform 1 0 4480 0 1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_28_32
timestamp 1698175906
transform 1 0 4928 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_28_34
timestamp 1698175906
transform 1 0 5152 0 1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_28_37
timestamp 1698175906
transform 1 0 5488 0 1 25088
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_28_45
timestamp 1698175906
transform 1 0 6384 0 1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_28_60
timestamp 1698175906
transform 1 0 8064 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_28_62
timestamp 1698175906
transform 1 0 8288 0 1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_28_121
timestamp 1698175906
transform 1 0 14896 0 1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_28_159
timestamp 1698175906
transform 1 0 19152 0 1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_28_177
timestamp 1698175906
transform 1 0 21168 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_28_228
timestamp 1698175906
transform 1 0 26880 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_28_232
timestamp 1698175906
transform 1 0 27328 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_28_234
timestamp 1698175906
transform 1 0 27552 0 1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_28_243
timestamp 1698175906
transform 1 0 28560 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_28_247
timestamp 1698175906
transform 1 0 29008 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_28_251
timestamp 1698175906
transform 1 0 29456 0 1 25088
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_28_317
timestamp 1698175906
transform 1 0 36848 0 1 25088
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_28_381
timestamp 1698175906
transform 1 0 44016 0 1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_28_387
timestamp 1698175906
transform 1 0 44688 0 1 25088
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_28_451
timestamp 1698175906
transform 1 0 51856 0 1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_28_457
timestamp 1698175906
transform 1 0 52528 0 1 25088
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_28_489
timestamp 1698175906
transform 1 0 56112 0 1 25088
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_28_505
timestamp 1698175906
transform 1 0 57904 0 1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_29_2
timestamp 1698175906
transform 1 0 1568 0 -1 26656
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_29_34
timestamp 1698175906
transform 1 0 5152 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_29_44
timestamp 1698175906
transform 1 0 6272 0 -1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_29_48
timestamp 1698175906
transform 1 0 6720 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_29_60
timestamp 1698175906
transform 1 0 8064 0 -1 26656
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_29_68
timestamp 1698175906
transform 1 0 8960 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_29_80
timestamp 1698175906
transform 1 0 10304 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_29_84
timestamp 1698175906
transform 1 0 10752 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_29_104
timestamp 1698175906
transform 1 0 12992 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_29_108
timestamp 1698175906
transform 1 0 13440 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_29_112
timestamp 1698175906
transform 1 0 13888 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_29_116
timestamp 1698175906
transform 1 0 14336 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_29_120
timestamp 1698175906
transform 1 0 14784 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_29_133
timestamp 1698175906
transform 1 0 16240 0 -1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_29_137
timestamp 1698175906
transform 1 0 16688 0 -1 26656
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_29_151
timestamp 1698175906
transform 1 0 18256 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_29_155
timestamp 1698175906
transform 1 0 18704 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_29_157
timestamp 1698175906
transform 1 0 18928 0 -1 26656
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_29_160
timestamp 1698175906
transform 1 0 19264 0 -1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_29_164
timestamp 1698175906
transform 1 0 19712 0 -1 26656
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_29_167
timestamp 1698175906
transform 1 0 20048 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_29_171
timestamp 1698175906
transform 1 0 20496 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_29_183
timestamp 1698175906
transform 1 0 21840 0 -1 26656
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_29_192
timestamp 1698175906
transform 1 0 22848 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_29_196
timestamp 1698175906
transform 1 0 23296 0 -1 26656
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_29_204
timestamp 1698175906
transform 1 0 24192 0 -1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_29_208
timestamp 1698175906
transform 1 0 24640 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_29_212
timestamp 1698175906
transform 1 0 25088 0 -1 26656
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_29_221
timestamp 1698175906
transform 1 0 26096 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_29_225
timestamp 1698175906
transform 1 0 26544 0 -1 26656
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_29_257
timestamp 1698175906
transform 1 0 30128 0 -1 26656
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_29_273
timestamp 1698175906
transform 1 0 31920 0 -1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_29_277
timestamp 1698175906
transform 1 0 32368 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_29_279
timestamp 1698175906
transform 1 0 32592 0 -1 26656
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_29_282
timestamp 1698175906
transform 1 0 32928 0 -1 26656
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_29_346
timestamp 1698175906
transform 1 0 40096 0 -1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_29_352
timestamp 1698175906
transform 1 0 40768 0 -1 26656
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_29_416
timestamp 1698175906
transform 1 0 47936 0 -1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_29_422
timestamp 1698175906
transform 1 0 48608 0 -1 26656
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_29_486
timestamp 1698175906
transform 1 0 55776 0 -1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_29_492
timestamp 1698175906
transform 1 0 56448 0 -1 26656
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_29_508
timestamp 1698175906
transform 1 0 58240 0 -1 26656
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_30_2
timestamp 1698175906
transform 1 0 1568 0 1 26656
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_30_18
timestamp 1698175906
transform 1 0 3360 0 1 26656
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_30_26
timestamp 1698175906
transform 1 0 4256 0 1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_30_32
timestamp 1698175906
transform 1 0 4928 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_30_34
timestamp 1698175906
transform 1 0 5152 0 1 26656
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_30_37
timestamp 1698175906
transform 1 0 5488 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_30_47
timestamp 1698175906
transform 1 0 6608 0 1 26656
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_30_63
timestamp 1698175906
transform 1 0 8400 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_30_65
timestamp 1698175906
transform 1 0 8624 0 1 26656
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_30_76
timestamp 1698175906
transform 1 0 9856 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_30_80
timestamp 1698175906
transform 1 0 10304 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_30_84
timestamp 1698175906
transform 1 0 10752 0 1 26656
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_30_92
timestamp 1698175906
transform 1 0 11648 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_30_94
timestamp 1698175906
transform 1 0 11872 0 1 26656
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_30_103
timestamp 1698175906
transform 1 0 12880 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_30_107
timestamp 1698175906
transform 1 0 13328 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_30_111
timestamp 1698175906
transform 1 0 13776 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_30_115
timestamp 1698175906
transform 1 0 14224 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_30_132
timestamp 1698175906
transform 1 0 16128 0 1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_30_138
timestamp 1698175906
transform 1 0 16800 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_30_142
timestamp 1698175906
transform 1 0 17248 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_30_146
timestamp 1698175906
transform 1 0 17696 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_30_158
timestamp 1698175906
transform 1 0 19040 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_30_162
timestamp 1698175906
transform 1 0 19488 0 1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_30_166
timestamp 1698175906
transform 1 0 19936 0 1 26656
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_30_169
timestamp 1698175906
transform 1 0 20272 0 1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_30_173
timestamp 1698175906
transform 1 0 20720 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_30_177
timestamp 1698175906
transform 1 0 21168 0 1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_30_181
timestamp 1698175906
transform 1 0 21616 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_30_185
timestamp 1698175906
transform 1 0 22064 0 1 26656
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_30_193
timestamp 1698175906
transform 1 0 22960 0 1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_30_197
timestamp 1698175906
transform 1 0 23408 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_30_199
timestamp 1698175906
transform 1 0 23632 0 1 26656
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_30_223
timestamp 1698175906
transform 1 0 26320 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_30_227
timestamp 1698175906
transform 1 0 26768 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_30_231
timestamp 1698175906
transform 1 0 27216 0 1 26656
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_30_239
timestamp 1698175906
transform 1 0 28112 0 1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_30_243
timestamp 1698175906
transform 1 0 28560 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_30_247
timestamp 1698175906
transform 1 0 29008 0 1 26656
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_30_311
timestamp 1698175906
transform 1 0 36176 0 1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_30_317
timestamp 1698175906
transform 1 0 36848 0 1 26656
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_30_381
timestamp 1698175906
transform 1 0 44016 0 1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_30_387
timestamp 1698175906
transform 1 0 44688 0 1 26656
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_30_451
timestamp 1698175906
transform 1 0 51856 0 1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_30_457
timestamp 1698175906
transform 1 0 52528 0 1 26656
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_30_489
timestamp 1698175906
transform 1 0 56112 0 1 26656
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_30_505
timestamp 1698175906
transform 1 0 57904 0 1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_31_8
timestamp 1698175906
transform 1 0 2240 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_31_12
timestamp 1698175906
transform 1 0 2688 0 -1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_31_16
timestamp 1698175906
transform 1 0 3136 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_31_27
timestamp 1698175906
transform 1 0 4368 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_31_29
timestamp 1698175906
transform 1 0 4592 0 -1 28224
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_31_86
timestamp 1698175906
transform 1 0 10976 0 -1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_31_90
timestamp 1698175906
transform 1 0 11424 0 -1 28224
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_31_142
timestamp 1698175906
transform 1 0 17248 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_31_144
timestamp 1698175906
transform 1 0 17472 0 -1 28224
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_31_182
timestamp 1698175906
transform 1 0 21728 0 -1 28224
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_31_192
timestamp 1698175906
transform 1 0 22848 0 -1 28224
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_31_220
timestamp 1698175906
transform 1 0 25984 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_31_222
timestamp 1698175906
transform 1 0 26208 0 -1 28224
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_31_237
timestamp 1698175906
transform 1 0 27888 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_31_241
timestamp 1698175906
transform 1 0 28336 0 -1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_31_245
timestamp 1698175906
transform 1 0 28784 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_31_263
timestamp 1698175906
transform 1 0 30800 0 -1 28224
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_31_279
timestamp 1698175906
transform 1 0 32592 0 -1 28224
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_31_282
timestamp 1698175906
transform 1 0 32928 0 -1 28224
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_31_346
timestamp 1698175906
transform 1 0 40096 0 -1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_31_352
timestamp 1698175906
transform 1 0 40768 0 -1 28224
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_31_416
timestamp 1698175906
transform 1 0 47936 0 -1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_31_422
timestamp 1698175906
transform 1 0 48608 0 -1 28224
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_31_486
timestamp 1698175906
transform 1 0 55776 0 -1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_31_492
timestamp 1698175906
transform 1 0 56448 0 -1 28224
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_31_508
timestamp 1698175906
transform 1 0 58240 0 -1 28224
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_32_2
timestamp 1698175906
transform 1 0 1568 0 1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_32_6
timestamp 1698175906
transform 1 0 2016 0 1 28224
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_32_25
timestamp 1698175906
transform 1 0 4144 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_32_29
timestamp 1698175906
transform 1 0 4592 0 1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_32_33
timestamp 1698175906
transform 1 0 5040 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_32_37
timestamp 1698175906
transform 1 0 5488 0 1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_32_41
timestamp 1698175906
transform 1 0 5936 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_32_91
timestamp 1698175906
transform 1 0 11536 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_32_95
timestamp 1698175906
transform 1 0 11984 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_32_99
timestamp 1698175906
transform 1 0 12432 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_32_103
timestamp 1698175906
transform 1 0 12880 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_32_107
timestamp 1698175906
transform 1 0 13328 0 1 28224
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_32_115
timestamp 1698175906
transform 1 0 14224 0 1 28224
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_32_127
timestamp 1698175906
transform 1 0 15568 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_32_139
timestamp 1698175906
transform 1 0 16912 0 1 28224
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_32_147
timestamp 1698175906
transform 1 0 17808 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_32_149
timestamp 1698175906
transform 1 0 18032 0 1 28224
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_32_157
timestamp 1698175906
transform 1 0 18928 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_32_161
timestamp 1698175906
transform 1 0 19376 0 1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_32_165
timestamp 1698175906
transform 1 0 19824 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_32_174
timestamp 1698175906
transform 1 0 20832 0 1 28224
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_32_190
timestamp 1698175906
transform 1 0 22624 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_32_210
timestamp 1698175906
transform 1 0 24864 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_32_214
timestamp 1698175906
transform 1 0 25312 0 1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_32_226
timestamp 1698175906
transform 1 0 26656 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_32_230
timestamp 1698175906
transform 1 0 27104 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_32_234
timestamp 1698175906
transform 1 0 27552 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_32_243
timestamp 1698175906
transform 1 0 28560 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_32_260
timestamp 1698175906
transform 1 0 30464 0 1 28224
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_32_292
timestamp 1698175906
transform 1 0 34048 0 1 28224
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_32_308
timestamp 1698175906
transform 1 0 35840 0 1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_32_312
timestamp 1698175906
transform 1 0 36288 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_32_314
timestamp 1698175906
transform 1 0 36512 0 1 28224
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_32_317
timestamp 1698175906
transform 1 0 36848 0 1 28224
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_32_381
timestamp 1698175906
transform 1 0 44016 0 1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_32_387
timestamp 1698175906
transform 1 0 44688 0 1 28224
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_32_451
timestamp 1698175906
transform 1 0 51856 0 1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_32_457
timestamp 1698175906
transform 1 0 52528 0 1 28224
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_32_489
timestamp 1698175906
transform 1 0 56112 0 1 28224
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_32_505
timestamp 1698175906
transform 1 0 57904 0 1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_33_2
timestamp 1698175906
transform 1 0 1568 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_33_6
timestamp 1698175906
transform 1 0 2016 0 -1 29792
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_33_47
timestamp 1698175906
transform 1 0 6608 0 -1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_33_68
timestamp 1698175906
transform 1 0 8960 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_33_88
timestamp 1698175906
transform 1 0 11200 0 -1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_33_102
timestamp 1698175906
transform 1 0 12768 0 -1 29792
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_33_114
timestamp 1698175906
transform 1 0 14112 0 -1 29792
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_33_125
timestamp 1698175906
transform 1 0 15344 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_33_129
timestamp 1698175906
transform 1 0 15792 0 -1 29792
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_33_137
timestamp 1698175906
transform 1 0 16688 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_33_139
timestamp 1698175906
transform 1 0 16912 0 -1 29792
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_33_142
timestamp 1698175906
transform 1 0 17248 0 -1 29792
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_33_150
timestamp 1698175906
transform 1 0 18144 0 -1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_33_154
timestamp 1698175906
transform 1 0 18592 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_33_156
timestamp 1698175906
transform 1 0 18816 0 -1 29792
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_33_159
timestamp 1698175906
transform 1 0 19152 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_33_172
timestamp 1698175906
transform 1 0 20608 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_33_182
timestamp 1698175906
transform 1 0 21728 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_33_186
timestamp 1698175906
transform 1 0 22176 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_33_190
timestamp 1698175906
transform 1 0 22624 0 -1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_33_194
timestamp 1698175906
transform 1 0 23072 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_33_196
timestamp 1698175906
transform 1 0 23296 0 -1 29792
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_33_199
timestamp 1698175906
transform 1 0 23632 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_33_208
timestamp 1698175906
transform 1 0 24640 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_33_212
timestamp 1698175906
transform 1 0 25088 0 -1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_33_216
timestamp 1698175906
transform 1 0 25536 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_33_220
timestamp 1698175906
transform 1 0 25984 0 -1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_33_224
timestamp 1698175906
transform 1 0 26432 0 -1 29792
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_33_227
timestamp 1698175906
transform 1 0 26768 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_33_255
timestamp 1698175906
transform 1 0 29904 0 -1 29792
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_33_271
timestamp 1698175906
transform 1 0 31696 0 -1 29792
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_33_279
timestamp 1698175906
transform 1 0 32592 0 -1 29792
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_33_282
timestamp 1698175906
transform 1 0 32928 0 -1 29792
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_33_290
timestamp 1698175906
transform 1 0 33824 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_33_292
timestamp 1698175906
transform 1 0 34048 0 -1 29792
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_33_330
timestamp 1698175906
transform 1 0 38304 0 -1 29792
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_33_346
timestamp 1698175906
transform 1 0 40096 0 -1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_33_352
timestamp 1698175906
transform 1 0 40768 0 -1 29792
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_33_416
timestamp 1698175906
transform 1 0 47936 0 -1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_33_422
timestamp 1698175906
transform 1 0 48608 0 -1 29792
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_33_486
timestamp 1698175906
transform 1 0 55776 0 -1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_33_492
timestamp 1698175906
transform 1 0 56448 0 -1 29792
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_33_508
timestamp 1698175906
transform 1 0 58240 0 -1 29792
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_34_14
timestamp 1698175906
transform 1 0 2912 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_34_18
timestamp 1698175906
transform 1 0 3360 0 1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_34_22
timestamp 1698175906
transform 1 0 3808 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_34_26
timestamp 1698175906
transform 1 0 4256 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_34_37
timestamp 1698175906
transform 1 0 5488 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_34_39
timestamp 1698175906
transform 1 0 5712 0 1 29792
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_34_51
timestamp 1698175906
transform 1 0 7056 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_34_53
timestamp 1698175906
transform 1 0 7280 0 1 29792
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_34_79
timestamp 1698175906
transform 1 0 10192 0 1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_34_85
timestamp 1698175906
transform 1 0 10864 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_34_98
timestamp 1698175906
transform 1 0 12320 0 1 29792
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_34_104
timestamp 1698175906
transform 1 0 12992 0 1 29792
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_34_107
timestamp 1698175906
transform 1 0 13328 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_34_111
timestamp 1698175906
transform 1 0 13776 0 1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_34_117
timestamp 1698175906
transform 1 0 14448 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_34_121
timestamp 1698175906
transform 1 0 14896 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_34_125
timestamp 1698175906
transform 1 0 15344 0 1 29792
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_34_186
timestamp 1698175906
transform 1 0 22176 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_34_221
timestamp 1698175906
transform 1 0 26096 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_34_225
timestamp 1698175906
transform 1 0 26544 0 1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_34_229
timestamp 1698175906
transform 1 0 26992 0 1 29792
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_34_232
timestamp 1698175906
transform 1 0 27328 0 1 29792
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_34_240
timestamp 1698175906
transform 1 0 28224 0 1 29792
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_34_243
timestamp 1698175906
transform 1 0 28560 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_34_247
timestamp 1698175906
transform 1 0 29008 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_34_251
timestamp 1698175906
transform 1 0 29456 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_34_253
timestamp 1698175906
transform 1 0 29680 0 1 29792
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_34_276
timestamp 1698175906
transform 1 0 32256 0 1 29792
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_34_292
timestamp 1698175906
transform 1 0 34048 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_34_294
timestamp 1698175906
transform 1 0 34272 0 1 29792
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_34_303
timestamp 1698175906
transform 1 0 35280 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_34_311
timestamp 1698175906
transform 1 0 36176 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_34_317
timestamp 1698175906
transform 1 0 36848 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_34_321
timestamp 1698175906
transform 1 0 37296 0 1 29792
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_34_387
timestamp 1698175906
transform 1 0 44688 0 1 29792
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_34_451
timestamp 1698175906
transform 1 0 51856 0 1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_34_457
timestamp 1698175906
transform 1 0 52528 0 1 29792
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_34_489
timestamp 1698175906
transform 1 0 56112 0 1 29792
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_34_505
timestamp 1698175906
transform 1 0 57904 0 1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_35_2
timestamp 1698175906
transform 1 0 1568 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_35_4
timestamp 1698175906
transform 1 0 1792 0 -1 31360
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_35_53
timestamp 1698175906
transform 1 0 7280 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_35_57
timestamp 1698175906
transform 1 0 7728 0 -1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_35_61
timestamp 1698175906
transform 1 0 8176 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_35_63
timestamp 1698175906
transform 1 0 8400 0 -1 31360
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_35_66
timestamp 1698175906
transform 1 0 8736 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_35_110
timestamp 1698175906
transform 1 0 13664 0 -1 31360
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_35_120
timestamp 1698175906
transform 1 0 14784 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_35_124
timestamp 1698175906
transform 1 0 15232 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_35_128
timestamp 1698175906
transform 1 0 15680 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_35_130
timestamp 1698175906
transform 1 0 15904 0 -1 31360
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_35_136
timestamp 1698175906
transform 1 0 16576 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_35_151
timestamp 1698175906
transform 1 0 18256 0 -1 31360
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_35_161
timestamp 1698175906
transform 1 0 19376 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_35_165
timestamp 1698175906
transform 1 0 19824 0 -1 31360
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_35_177
timestamp 1698175906
transform 1 0 21168 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_35_181
timestamp 1698175906
transform 1 0 21616 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_35_185
timestamp 1698175906
transform 1 0 22064 0 -1 31360
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_35_228
timestamp 1698175906
transform 1 0 26880 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_35_240
timestamp 1698175906
transform 1 0 28224 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_35_242
timestamp 1698175906
transform 1 0 28448 0 -1 31360
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_35_251
timestamp 1698175906
transform 1 0 29456 0 -1 31360
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_35_267
timestamp 1698175906
transform 1 0 31248 0 -1 31360
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_35_275
timestamp 1698175906
transform 1 0 32144 0 -1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_35_279
timestamp 1698175906
transform 1 0 32592 0 -1 31360
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_35_333
timestamp 1698175906
transform 1 0 38640 0 -1 31360
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_35_349
timestamp 1698175906
transform 1 0 40432 0 -1 31360
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_35_352
timestamp 1698175906
transform 1 0 40768 0 -1 31360
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_35_416
timestamp 1698175906
transform 1 0 47936 0 -1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_35_422
timestamp 1698175906
transform 1 0 48608 0 -1 31360
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_35_486
timestamp 1698175906
transform 1 0 55776 0 -1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_35_492
timestamp 1698175906
transform 1 0 56448 0 -1 31360
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_35_508
timestamp 1698175906
transform 1 0 58240 0 -1 31360
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_36_2
timestamp 1698175906
transform 1 0 1568 0 1 31360
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_36_10
timestamp 1698175906
transform 1 0 2464 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_36_28
timestamp 1698175906
transform 1 0 4480 0 1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_36_32
timestamp 1698175906
transform 1 0 4928 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_36_34
timestamp 1698175906
transform 1 0 5152 0 1 31360
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_36_37
timestamp 1698175906
transform 1 0 5488 0 1 31360
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_36_53
timestamp 1698175906
transform 1 0 7280 0 1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_36_57
timestamp 1698175906
transform 1 0 7728 0 1 31360
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_36_115
timestamp 1698175906
transform 1 0 14224 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_36_126
timestamp 1698175906
transform 1 0 15456 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_36_160
timestamp 1698175906
transform 1 0 19264 0 1 31360
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_36_177
timestamp 1698175906
transform 1 0 21168 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_36_181
timestamp 1698175906
transform 1 0 21616 0 1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_36_185
timestamp 1698175906
transform 1 0 22064 0 1 31360
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_36_194
timestamp 1698175906
transform 1 0 23072 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_36_243
timestamp 1698175906
transform 1 0 28560 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_36_255
timestamp 1698175906
transform 1 0 29904 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_36_257
timestamp 1698175906
transform 1 0 30128 0 1 31360
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_36_266
timestamp 1698175906
transform 1 0 31136 0 1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_36_270
timestamp 1698175906
transform 1 0 31584 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_36_272
timestamp 1698175906
transform 1 0 31808 0 1 31360
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_36_310
timestamp 1698175906
transform 1 0 36064 0 1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_36_314
timestamp 1698175906
transform 1 0 36512 0 1 31360
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_36_354
timestamp 1698175906
transform 1 0 40992 0 1 31360
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_36_370
timestamp 1698175906
transform 1 0 42784 0 1 31360
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_36_378
timestamp 1698175906
transform 1 0 43680 0 1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_36_382
timestamp 1698175906
transform 1 0 44128 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_36_384
timestamp 1698175906
transform 1 0 44352 0 1 31360
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_36_387
timestamp 1698175906
transform 1 0 44688 0 1 31360
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_36_451
timestamp 1698175906
transform 1 0 51856 0 1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_36_457
timestamp 1698175906
transform 1 0 52528 0 1 31360
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_36_489
timestamp 1698175906
transform 1 0 56112 0 1 31360
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_36_505
timestamp 1698175906
transform 1 0 57904 0 1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_37_2
timestamp 1698175906
transform 1 0 1568 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_37_51
timestamp 1698175906
transform 1 0 7056 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_37_55
timestamp 1698175906
transform 1 0 7504 0 -1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_37_59
timestamp 1698175906
transform 1 0 7952 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_37_61
timestamp 1698175906
transform 1 0 8176 0 -1 32928
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_37_72
timestamp 1698175906
transform 1 0 9408 0 -1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_37_76
timestamp 1698175906
transform 1 0 9856 0 -1 32928
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_37_110
timestamp 1698175906
transform 1 0 13664 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_37_122
timestamp 1698175906
transform 1 0 15008 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_37_126
timestamp 1698175906
transform 1 0 15456 0 -1 32928
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_37_136
timestamp 1698175906
transform 1 0 16576 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_37_157
timestamp 1698175906
transform 1 0 18928 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_37_161
timestamp 1698175906
transform 1 0 19376 0 -1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_37_167
timestamp 1698175906
transform 1 0 20048 0 -1 32928
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_37_175
timestamp 1698175906
transform 1 0 20944 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_37_177
timestamp 1698175906
transform 1 0 21168 0 -1 32928
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_37_203
timestamp 1698175906
transform 1 0 24080 0 -1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_37_207
timestamp 1698175906
transform 1 0 24528 0 -1 32928
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_37_244
timestamp 1698175906
transform 1 0 28672 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_37_248
timestamp 1698175906
transform 1 0 29120 0 -1 32928
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_37_347
timestamp 1698175906
transform 1 0 40208 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_37_349
timestamp 1698175906
transform 1 0 40432 0 -1 32928
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_37_360
timestamp 1698175906
transform 1 0 41664 0 -1 32928
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_37_392
timestamp 1698175906
transform 1 0 45248 0 -1 32928
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_37_408
timestamp 1698175906
transform 1 0 47040 0 -1 32928
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_37_416
timestamp 1698175906
transform 1 0 47936 0 -1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_37_422
timestamp 1698175906
transform 1 0 48608 0 -1 32928
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_37_486
timestamp 1698175906
transform 1 0 55776 0 -1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_37_492
timestamp 1698175906
transform 1 0 56448 0 -1 32928
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_37_508
timestamp 1698175906
transform 1 0 58240 0 -1 32928
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_38_8
timestamp 1698175906
transform 1 0 2240 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_38_23
timestamp 1698175906
transform 1 0 3920 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_38_37
timestamp 1698175906
transform 1 0 5488 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_38_39
timestamp 1698175906
transform 1 0 5712 0 1 32928
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_38_72
timestamp 1698175906
transform 1 0 9408 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_38_76
timestamp 1698175906
transform 1 0 9856 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_38_80
timestamp 1698175906
transform 1 0 10304 0 1 32928
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_38_88
timestamp 1698175906
transform 1 0 11200 0 1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_38_92
timestamp 1698175906
transform 1 0 11648 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_38_94
timestamp 1698175906
transform 1 0 11872 0 1 32928
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_38_97
timestamp 1698175906
transform 1 0 12208 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_38_101
timestamp 1698175906
transform 1 0 12656 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_38_107
timestamp 1698175906
transform 1 0 13328 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_38_109
timestamp 1698175906
transform 1 0 13552 0 1 32928
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_38_112
timestamp 1698175906
transform 1 0 13888 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_38_116
timestamp 1698175906
transform 1 0 14336 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_38_120
timestamp 1698175906
transform 1 0 14784 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_38_124
timestamp 1698175906
transform 1 0 15232 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_38_128
timestamp 1698175906
transform 1 0 15680 0 1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_38_132
timestamp 1698175906
transform 1 0 16128 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_38_136
timestamp 1698175906
transform 1 0 16576 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_38_138
timestamp 1698175906
transform 1 0 16800 0 1 32928
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_38_160
timestamp 1698175906
transform 1 0 19264 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_38_164
timestamp 1698175906
transform 1 0 19712 0 1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_38_168
timestamp 1698175906
transform 1 0 20160 0 1 32928
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_38_171
timestamp 1698175906
transform 1 0 20496 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_38_177
timestamp 1698175906
transform 1 0 21168 0 1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_38_183
timestamp 1698175906
transform 1 0 21840 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_38_187
timestamp 1698175906
transform 1 0 22288 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_38_231
timestamp 1698175906
transform 1 0 27216 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_38_242
timestamp 1698175906
transform 1 0 28448 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_38_244
timestamp 1698175906
transform 1 0 28672 0 1 32928
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_38_247
timestamp 1698175906
transform 1 0 29008 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_38_251
timestamp 1698175906
transform 1 0 29456 0 1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_38_255
timestamp 1698175906
transform 1 0 29904 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_38_265
timestamp 1698175906
transform 1 0 31024 0 1 32928
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_38_305
timestamp 1698175906
transform 1 0 35504 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_38_317
timestamp 1698175906
transform 1 0 36848 0 1 32928
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_38_359
timestamp 1698175906
transform 1 0 41552 0 1 32928
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_38_375
timestamp 1698175906
transform 1 0 43344 0 1 32928
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_38_383
timestamp 1698175906
transform 1 0 44240 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_38_387
timestamp 1698175906
transform 1 0 44688 0 1 32928
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_38_451
timestamp 1698175906
transform 1 0 51856 0 1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_38_457
timestamp 1698175906
transform 1 0 52528 0 1 32928
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_38_489
timestamp 1698175906
transform 1 0 56112 0 1 32928
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_38_505
timestamp 1698175906
transform 1 0 57904 0 1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_39_8
timestamp 1698175906
transform 1 0 2240 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_39_12
timestamp 1698175906
transform 1 0 2688 0 -1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_39_24
timestamp 1698175906
transform 1 0 4032 0 -1 34496
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_39_32
timestamp 1698175906
transform 1 0 4928 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_39_34
timestamp 1698175906
transform 1 0 5152 0 -1 34496
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_39_43
timestamp 1698175906
transform 1 0 6160 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_39_45
timestamp 1698175906
transform 1 0 6384 0 -1 34496
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_39_48
timestamp 1698175906
transform 1 0 6720 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_39_60
timestamp 1698175906
transform 1 0 8064 0 -1 34496
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_39_69
timestamp 1698175906
transform 1 0 9072 0 -1 34496
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_39_85
timestamp 1698175906
transform 1 0 10864 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_39_89
timestamp 1698175906
transform 1 0 11312 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_39_101
timestamp 1698175906
transform 1 0 12656 0 -1 34496
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_39_134
timestamp 1698175906
transform 1 0 16352 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_39_138
timestamp 1698175906
transform 1 0 16800 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_39_147
timestamp 1698175906
transform 1 0 17808 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_39_159
timestamp 1698175906
transform 1 0 19152 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_39_161
timestamp 1698175906
transform 1 0 19376 0 -1 34496
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_39_205
timestamp 1698175906
transform 1 0 24304 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_39_207
timestamp 1698175906
transform 1 0 24528 0 -1 34496
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_39_227
timestamp 1698175906
transform 1 0 26768 0 -1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_39_243
timestamp 1698175906
transform 1 0 28560 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_39_247
timestamp 1698175906
transform 1 0 29008 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_39_251
timestamp 1698175906
transform 1 0 29456 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_39_255
timestamp 1698175906
transform 1 0 29904 0 -1 34496
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_39_264
timestamp 1698175906
transform 1 0 30912 0 -1 34496
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_39_322
timestamp 1698175906
transform 1 0 37408 0 -1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_39_326
timestamp 1698175906
transform 1 0 37856 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_39_328
timestamp 1698175906
transform 1 0 38080 0 -1 34496
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_39_343
timestamp 1698175906
transform 1 0 39760 0 -1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_39_347
timestamp 1698175906
transform 1 0 40208 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_39_349
timestamp 1698175906
transform 1 0 40432 0 -1 34496
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_39_352
timestamp 1698175906
transform 1 0 40768 0 -1 34496
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_39_416
timestamp 1698175906
transform 1 0 47936 0 -1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_39_422
timestamp 1698175906
transform 1 0 48608 0 -1 34496
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_39_486
timestamp 1698175906
transform 1 0 55776 0 -1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_39_492
timestamp 1698175906
transform 1 0 56448 0 -1 34496
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_39_508
timestamp 1698175906
transform 1 0 58240 0 -1 34496
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_40_2
timestamp 1698175906
transform 1 0 1568 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_40_6
timestamp 1698175906
transform 1 0 2016 0 1 34496
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_40_16
timestamp 1698175906
transform 1 0 3136 0 1 34496
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_40_32
timestamp 1698175906
transform 1 0 4928 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_40_34
timestamp 1698175906
transform 1 0 5152 0 1 34496
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_40_67
timestamp 1698175906
transform 1 0 8848 0 1 34496
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_40_93
timestamp 1698175906
transform 1 0 11760 0 1 34496
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_40_101
timestamp 1698175906
transform 1 0 12656 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_40_164
timestamp 1698175906
transform 1 0 19712 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_40_166
timestamp 1698175906
transform 1 0 19936 0 1 34496
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_40_177
timestamp 1698175906
transform 1 0 21168 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_40_179
timestamp 1698175906
transform 1 0 21392 0 1 34496
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_40_241
timestamp 1698175906
transform 1 0 28336 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_40_247
timestamp 1698175906
transform 1 0 29008 0 1 34496
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_40_266
timestamp 1698175906
transform 1 0 31136 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_40_268
timestamp 1698175906
transform 1 0 31360 0 1 34496
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_40_295
timestamp 1698175906
transform 1 0 34384 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_40_354
timestamp 1698175906
transform 1 0 40992 0 1 34496
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_40_370
timestamp 1698175906
transform 1 0 42784 0 1 34496
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_40_378
timestamp 1698175906
transform 1 0 43680 0 1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_40_382
timestamp 1698175906
transform 1 0 44128 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_40_384
timestamp 1698175906
transform 1 0 44352 0 1 34496
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_40_387
timestamp 1698175906
transform 1 0 44688 0 1 34496
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_40_451
timestamp 1698175906
transform 1 0 51856 0 1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_40_457
timestamp 1698175906
transform 1 0 52528 0 1 34496
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_40_489
timestamp 1698175906
transform 1 0 56112 0 1 34496
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_40_505
timestamp 1698175906
transform 1 0 57904 0 1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_41_2
timestamp 1698175906
transform 1 0 1568 0 -1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_41_6
timestamp 1698175906
transform 1 0 2016 0 -1 36064
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_41_23
timestamp 1698175906
transform 1 0 3920 0 -1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_41_27
timestamp 1698175906
transform 1 0 4368 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_41_31
timestamp 1698175906
transform 1 0 4816 0 -1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_41_35
timestamp 1698175906
transform 1 0 5264 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_41_37
timestamp 1698175906
transform 1 0 5488 0 -1 36064
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_41_46
timestamp 1698175906
transform 1 0 6496 0 -1 36064
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_41_54
timestamp 1698175906
transform 1 0 7392 0 -1 36064
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_41_63
timestamp 1698175906
transform 1 0 8400 0 -1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_41_67
timestamp 1698175906
transform 1 0 8848 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_41_69
timestamp 1698175906
transform 1 0 9072 0 -1 36064
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_41_72
timestamp 1698175906
transform 1 0 9408 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_41_74
timestamp 1698175906
transform 1 0 9632 0 -1 36064
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_41_82
timestamp 1698175906
transform 1 0 10528 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_41_86
timestamp 1698175906
transform 1 0 10976 0 -1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_41_92
timestamp 1698175906
transform 1 0 11648 0 -1 36064
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_41_98
timestamp 1698175906
transform 1 0 12320 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_41_102
timestamp 1698175906
transform 1 0 12768 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_41_106
timestamp 1698175906
transform 1 0 13216 0 -1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_41_123
timestamp 1698175906
transform 1 0 15120 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_41_127
timestamp 1698175906
transform 1 0 15568 0 -1 36064
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_41_135
timestamp 1698175906
transform 1 0 16464 0 -1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_41_139
timestamp 1698175906
transform 1 0 16912 0 -1 36064
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_41_142
timestamp 1698175906
transform 1 0 17248 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_41_162
timestamp 1698175906
transform 1 0 19488 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_41_221
timestamp 1698175906
transform 1 0 26096 0 -1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_41_225
timestamp 1698175906
transform 1 0 26544 0 -1 36064
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_41_228
timestamp 1698175906
transform 1 0 26880 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_41_243
timestamp 1698175906
transform 1 0 28560 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_41_247
timestamp 1698175906
transform 1 0 29008 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_41_251
timestamp 1698175906
transform 1 0 29456 0 -1 36064
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_41_267
timestamp 1698175906
transform 1 0 31248 0 -1 36064
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_41_275
timestamp 1698175906
transform 1 0 32144 0 -1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_41_279
timestamp 1698175906
transform 1 0 32592 0 -1 36064
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_41_282
timestamp 1698175906
transform 1 0 32928 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_41_345
timestamp 1698175906
transform 1 0 39984 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_41_347
timestamp 1698175906
transform 1 0 40208 0 -1 36064
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_41_360
timestamp 1698175906
transform 1 0 41664 0 -1 36064
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_41_392
timestamp 1698175906
transform 1 0 45248 0 -1 36064
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_41_408
timestamp 1698175906
transform 1 0 47040 0 -1 36064
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_41_416
timestamp 1698175906
transform 1 0 47936 0 -1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_41_422
timestamp 1698175906
transform 1 0 48608 0 -1 36064
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_41_486
timestamp 1698175906
transform 1 0 55776 0 -1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_41_492
timestamp 1698175906
transform 1 0 56448 0 -1 36064
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_41_508
timestamp 1698175906
transform 1 0 58240 0 -1 36064
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_42_2
timestamp 1698175906
transform 1 0 1568 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_42_29
timestamp 1698175906
transform 1 0 4592 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_42_33
timestamp 1698175906
transform 1 0 5040 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_42_43
timestamp 1698175906
transform 1 0 6160 0 1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_42_66
timestamp 1698175906
transform 1 0 8736 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_42_70
timestamp 1698175906
transform 1 0 9184 0 1 36064
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_42_78
timestamp 1698175906
transform 1 0 10080 0 1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_42_84
timestamp 1698175906
transform 1 0 10752 0 1 36064
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_42_100
timestamp 1698175906
transform 1 0 12544 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_42_102
timestamp 1698175906
transform 1 0 12768 0 1 36064
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_42_107
timestamp 1698175906
transform 1 0 13328 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_42_109
timestamp 1698175906
transform 1 0 13552 0 1 36064
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_42_117
timestamp 1698175906
transform 1 0 14448 0 1 36064
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_42_133
timestamp 1698175906
transform 1 0 16240 0 1 36064
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_42_141
timestamp 1698175906
transform 1 0 17136 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_42_143
timestamp 1698175906
transform 1 0 17360 0 1 36064
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_42_153
timestamp 1698175906
transform 1 0 18480 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_42_155
timestamp 1698175906
transform 1 0 18704 0 1 36064
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_42_158
timestamp 1698175906
transform 1 0 19040 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_42_162
timestamp 1698175906
transform 1 0 19488 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_42_166
timestamp 1698175906
transform 1 0 19936 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_42_177
timestamp 1698175906
transform 1 0 21168 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_42_181
timestamp 1698175906
transform 1 0 21616 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_42_232
timestamp 1698175906
transform 1 0 27328 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_42_236
timestamp 1698175906
transform 1 0 27776 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_42_247
timestamp 1698175906
transform 1 0 29008 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_42_251
timestamp 1698175906
transform 1 0 29456 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_42_255
timestamp 1698175906
transform 1 0 29904 0 1 36064
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_42_263
timestamp 1698175906
transform 1 0 30800 0 1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_42_267
timestamp 1698175906
transform 1 0 31248 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_42_269
timestamp 1698175906
transform 1 0 31472 0 1 36064
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_42_278
timestamp 1698175906
transform 1 0 32480 0 1 36064
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_42_313
timestamp 1698175906
transform 1 0 36400 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_42_355
timestamp 1698175906
transform 1 0 41104 0 1 36064
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_42_371
timestamp 1698175906
transform 1 0 42896 0 1 36064
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_42_379
timestamp 1698175906
transform 1 0 43792 0 1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_42_383
timestamp 1698175906
transform 1 0 44240 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_42_387
timestamp 1698175906
transform 1 0 44688 0 1 36064
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_42_451
timestamp 1698175906
transform 1 0 51856 0 1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_42_457
timestamp 1698175906
transform 1 0 52528 0 1 36064
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_42_489
timestamp 1698175906
transform 1 0 56112 0 1 36064
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_42_505
timestamp 1698175906
transform 1 0 57904 0 1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_43_8
timestamp 1698175906
transform 1 0 2240 0 -1 37632
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_43_14
timestamp 1698175906
transform 1 0 2912 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_43_18
timestamp 1698175906
transform 1 0 3360 0 -1 37632
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_43_34
timestamp 1698175906
transform 1 0 5152 0 -1 37632
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_43_42
timestamp 1698175906
transform 1 0 6048 0 -1 37632
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_43_45
timestamp 1698175906
transform 1 0 6384 0 -1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_43_49
timestamp 1698175906
transform 1 0 6832 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_43_51
timestamp 1698175906
transform 1 0 7056 0 -1 37632
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_43_83
timestamp 1698175906
transform 1 0 10640 0 -1 37632
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_43_91
timestamp 1698175906
transform 1 0 11536 0 -1 37632
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_43_98
timestamp 1698175906
transform 1 0 12320 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_43_102
timestamp 1698175906
transform 1 0 12768 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_43_106
timestamp 1698175906
transform 1 0 13216 0 -1 37632
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_43_114
timestamp 1698175906
transform 1 0 14112 0 -1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_43_118
timestamp 1698175906
transform 1 0 14560 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_43_137
timestamp 1698175906
transform 1 0 16688 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_43_139
timestamp 1698175906
transform 1 0 16912 0 -1 37632
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_43_142
timestamp 1698175906
transform 1 0 17248 0 -1 37632
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_43_149
timestamp 1698175906
transform 1 0 18032 0 -1 37632
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_43_155
timestamp 1698175906
transform 1 0 18704 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_43_162
timestamp 1698175906
transform 1 0 19488 0 -1 37632
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_43_212
timestamp 1698175906
transform 1 0 25088 0 -1 37632
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_43_239
timestamp 1698175906
transform 1 0 28112 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_43_243
timestamp 1698175906
transform 1 0 28560 0 -1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_43_278
timestamp 1698175906
transform 1 0 32480 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_43_282
timestamp 1698175906
transform 1 0 32928 0 -1 37632
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_43_290
timestamp 1698175906
transform 1 0 33824 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_43_339
timestamp 1698175906
transform 1 0 39312 0 -1 37632
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_43_352
timestamp 1698175906
transform 1 0 40768 0 -1 37632
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_43_416
timestamp 1698175906
transform 1 0 47936 0 -1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_43_422
timestamp 1698175906
transform 1 0 48608 0 -1 37632
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_43_486
timestamp 1698175906
transform 1 0 55776 0 -1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_43_492
timestamp 1698175906
transform 1 0 56448 0 -1 37632
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_43_508
timestamp 1698175906
transform 1 0 58240 0 -1 37632
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_44_8
timestamp 1698175906
transform 1 0 2240 0 1 37632
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_44_33
timestamp 1698175906
transform 1 0 5040 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_44_62
timestamp 1698175906
transform 1 0 8288 0 1 37632
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_44_80
timestamp 1698175906
transform 1 0 10304 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_44_100
timestamp 1698175906
transform 1 0 12544 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_44_104
timestamp 1698175906
transform 1 0 12992 0 1 37632
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_44_132
timestamp 1698175906
transform 1 0 16128 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_44_136
timestamp 1698175906
transform 1 0 16576 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_44_138
timestamp 1698175906
transform 1 0 16800 0 1 37632
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_44_148
timestamp 1698175906
transform 1 0 17920 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_44_160
timestamp 1698175906
transform 1 0 19264 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_44_173
timestamp 1698175906
transform 1 0 20720 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_44_177
timestamp 1698175906
transform 1 0 21168 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_44_179
timestamp 1698175906
transform 1 0 21392 0 1 37632
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_44_182
timestamp 1698175906
transform 1 0 21728 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_44_186
timestamp 1698175906
transform 1 0 22176 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_44_190
timestamp 1698175906
transform 1 0 22624 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_44_194
timestamp 1698175906
transform 1 0 23072 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_44_198
timestamp 1698175906
transform 1 0 23520 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_44_247
timestamp 1698175906
transform 1 0 29008 0 1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_44_251
timestamp 1698175906
transform 1 0 29456 0 1 37632
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_44_263
timestamp 1698175906
transform 1 0 30800 0 1 37632
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_44_271
timestamp 1698175906
transform 1 0 31696 0 1 37632
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_44_277
timestamp 1698175906
transform 1 0 32368 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_44_279
timestamp 1698175906
transform 1 0 32592 0 1 37632
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_44_296
timestamp 1698175906
transform 1 0 34496 0 1 37632
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_44_312
timestamp 1698175906
transform 1 0 36288 0 1 37632
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_44_317
timestamp 1698175906
transform 1 0 36848 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_44_333
timestamp 1698175906
transform 1 0 38640 0 1 37632
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_44_365
timestamp 1698175906
transform 1 0 42224 0 1 37632
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_44_381
timestamp 1698175906
transform 1 0 44016 0 1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_44_387
timestamp 1698175906
transform 1 0 44688 0 1 37632
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_44_451
timestamp 1698175906
transform 1 0 51856 0 1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_44_457
timestamp 1698175906
transform 1 0 52528 0 1 37632
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_44_489
timestamp 1698175906
transform 1 0 56112 0 1 37632
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_44_505
timestamp 1698175906
transform 1 0 57904 0 1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_45_2
timestamp 1698175906
transform 1 0 1568 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_45_6
timestamp 1698175906
transform 1 0 2016 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_45_14
timestamp 1698175906
transform 1 0 2912 0 -1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_45_24
timestamp 1698175906
transform 1 0 4032 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_45_28
timestamp 1698175906
transform 1 0 4480 0 -1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_45_32
timestamp 1698175906
transform 1 0 4928 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_45_34
timestamp 1698175906
transform 1 0 5152 0 -1 39200
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_45_63
timestamp 1698175906
transform 1 0 8400 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_45_67
timestamp 1698175906
transform 1 0 8848 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_45_69
timestamp 1698175906
transform 1 0 9072 0 -1 39200
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_45_72
timestamp 1698175906
transform 1 0 9408 0 -1 39200
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_45_88
timestamp 1698175906
transform 1 0 11200 0 -1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_45_106
timestamp 1698175906
transform 1 0 13216 0 -1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_45_110
timestamp 1698175906
transform 1 0 13664 0 -1 39200
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_45_128
timestamp 1698175906
transform 1 0 15680 0 -1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_45_134
timestamp 1698175906
transform 1 0 16352 0 -1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_45_138
timestamp 1698175906
transform 1 0 16800 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_45_142
timestamp 1698175906
transform 1 0 17248 0 -1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_45_146
timestamp 1698175906
transform 1 0 17696 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_45_150
timestamp 1698175906
transform 1 0 18144 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_45_152
timestamp 1698175906
transform 1 0 18368 0 -1 39200
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_45_155
timestamp 1698175906
transform 1 0 18704 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_45_159
timestamp 1698175906
transform 1 0 19152 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_45_163
timestamp 1698175906
transform 1 0 19600 0 -1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_45_167
timestamp 1698175906
transform 1 0 20048 0 -1 39200
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_45_170
timestamp 1698175906
transform 1 0 20384 0 -1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_45_193
timestamp 1698175906
transform 1 0 22960 0 -1 39200
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_45_202
timestamp 1698175906
transform 1 0 23968 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_45_206
timestamp 1698175906
transform 1 0 24416 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_45_235
timestamp 1698175906
transform 1 0 27664 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_45_239
timestamp 1698175906
transform 1 0 28112 0 -1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_45_243
timestamp 1698175906
transform 1 0 28560 0 -1 39200
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_45_246
timestamp 1698175906
transform 1 0 28896 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_45_250
timestamp 1698175906
transform 1 0 29344 0 -1 39200
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_45_258
timestamp 1698175906
transform 1 0 30240 0 -1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_45_262
timestamp 1698175906
transform 1 0 30688 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_45_282
timestamp 1698175906
transform 1 0 32928 0 -1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_45_318
timestamp 1698175906
transform 1 0 36960 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_45_320
timestamp 1698175906
transform 1 0 37184 0 -1 39200
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_45_352
timestamp 1698175906
transform 1 0 40768 0 -1 39200
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_45_416
timestamp 1698175906
transform 1 0 47936 0 -1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_45_422
timestamp 1698175906
transform 1 0 48608 0 -1 39200
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_45_486
timestamp 1698175906
transform 1 0 55776 0 -1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_45_492
timestamp 1698175906
transform 1 0 56448 0 -1 39200
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_45_508
timestamp 1698175906
transform 1 0 58240 0 -1 39200
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_46_2
timestamp 1698175906
transform 1 0 1568 0 1 39200
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_46_10
timestamp 1698175906
transform 1 0 2464 0 1 39200
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_46_37
timestamp 1698175906
transform 1 0 5488 0 1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_46_41
timestamp 1698175906
transform 1 0 5936 0 1 39200
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_46_76
timestamp 1698175906
transform 1 0 9856 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_46_92
timestamp 1698175906
transform 1 0 11648 0 1 39200
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_46_100
timestamp 1698175906
transform 1 0 12544 0 1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_46_104
timestamp 1698175906
transform 1 0 12992 0 1 39200
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_46_107
timestamp 1698175906
transform 1 0 13328 0 1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_46_111
timestamp 1698175906
transform 1 0 13776 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_46_113
timestamp 1698175906
transform 1 0 14000 0 1 39200
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_46_116
timestamp 1698175906
transform 1 0 14336 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_46_160
timestamp 1698175906
transform 1 0 19264 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_46_164
timestamp 1698175906
transform 1 0 19712 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_46_168
timestamp 1698175906
transform 1 0 20160 0 1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_46_172
timestamp 1698175906
transform 1 0 20608 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_46_174
timestamp 1698175906
transform 1 0 20832 0 1 39200
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_46_191
timestamp 1698175906
transform 1 0 22736 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_46_232
timestamp 1698175906
transform 1 0 27328 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_46_244
timestamp 1698175906
transform 1 0 28672 0 1 39200
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_46_247
timestamp 1698175906
transform 1 0 29008 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_46_249
timestamp 1698175906
transform 1 0 29232 0 1 39200
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_46_307
timestamp 1698175906
transform 1 0 35728 0 1 39200
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_46_317
timestamp 1698175906
transform 1 0 36848 0 1 39200
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_46_381
timestamp 1698175906
transform 1 0 44016 0 1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_46_387
timestamp 1698175906
transform 1 0 44688 0 1 39200
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_46_451
timestamp 1698175906
transform 1 0 51856 0 1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_46_457
timestamp 1698175906
transform 1 0 52528 0 1 39200
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_46_489
timestamp 1698175906
transform 1 0 56112 0 1 39200
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_46_505
timestamp 1698175906
transform 1 0 57904 0 1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_47_8
timestamp 1698175906
transform 1 0 2240 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_47_12
timestamp 1698175906
transform 1 0 2688 0 -1 40768
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_47_16
timestamp 1698175906
transform 1 0 3136 0 -1 40768
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_47_72
timestamp 1698175906
transform 1 0 9408 0 -1 40768
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_47_109
timestamp 1698175906
transform 1 0 13552 0 -1 40768
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_47_113
timestamp 1698175906
transform 1 0 14000 0 -1 40768
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_47_122
timestamp 1698175906
transform 1 0 15008 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_47_139
timestamp 1698175906
transform 1 0 16912 0 -1 40768
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_47_148
timestamp 1698175906
transform 1 0 17920 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_47_163
timestamp 1698175906
transform 1 0 19600 0 -1 40768
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_47_171
timestamp 1698175906
transform 1 0 20496 0 -1 40768
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_47_177
timestamp 1698175906
transform 1 0 21168 0 -1 40768
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_47_185
timestamp 1698175906
transform 1 0 22064 0 -1 40768
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_47_191
timestamp 1698175906
transform 1 0 22736 0 -1 40768
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_47_199
timestamp 1698175906
transform 1 0 23632 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_47_201
timestamp 1698175906
transform 1 0 23856 0 -1 40768
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_47_204
timestamp 1698175906
transform 1 0 24192 0 -1 40768
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_47_208
timestamp 1698175906
transform 1 0 24640 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_47_228
timestamp 1698175906
transform 1 0 26880 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_47_230
timestamp 1698175906
transform 1 0 27104 0 -1 40768
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_47_233
timestamp 1698175906
transform 1 0 27440 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_47_282
timestamp 1698175906
transform 1 0 32928 0 -1 40768
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_47_290
timestamp 1698175906
transform 1 0 33824 0 -1 40768
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_47_309
timestamp 1698175906
transform 1 0 35952 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_47_313
timestamp 1698175906
transform 1 0 36400 0 -1 40768
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_47_346
timestamp 1698175906
transform 1 0 40096 0 -1 40768
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_47_352
timestamp 1698175906
transform 1 0 40768 0 -1 40768
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_47_416
timestamp 1698175906
transform 1 0 47936 0 -1 40768
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_47_422
timestamp 1698175906
transform 1 0 48608 0 -1 40768
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_47_486
timestamp 1698175906
transform 1 0 55776 0 -1 40768
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_47_492
timestamp 1698175906
transform 1 0 56448 0 -1 40768
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_47_508
timestamp 1698175906
transform 1 0 58240 0 -1 40768
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_48_14
timestamp 1698175906
transform 1 0 2912 0 1 40768
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_48_30
timestamp 1698175906
transform 1 0 4704 0 1 40768
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_48_34
timestamp 1698175906
transform 1 0 5152 0 1 40768
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_48_37
timestamp 1698175906
transform 1 0 5488 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_48_87
timestamp 1698175906
transform 1 0 11088 0 1 40768
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_48_91
timestamp 1698175906
transform 1 0 11536 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_48_102
timestamp 1698175906
transform 1 0 12768 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_48_104
timestamp 1698175906
transform 1 0 12992 0 1 40768
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_48_107
timestamp 1698175906
transform 1 0 13328 0 1 40768
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_48_120
timestamp 1698175906
transform 1 0 14784 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_48_124
timestamp 1698175906
transform 1 0 15232 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_48_168
timestamp 1698175906
transform 1 0 20160 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_48_187
timestamp 1698175906
transform 1 0 22288 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_48_191
timestamp 1698175906
transform 1 0 22736 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_48_257
timestamp 1698175906
transform 1 0 30128 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_48_261
timestamp 1698175906
transform 1 0 30576 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_48_263
timestamp 1698175906
transform 1 0 30800 0 1 40768
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_48_296
timestamp 1698175906
transform 1 0 34496 0 1 40768
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_48_313
timestamp 1698175906
transform 1 0 36400 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_48_317
timestamp 1698175906
transform 1 0 36848 0 1 40768
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_48_381
timestamp 1698175906
transform 1 0 44016 0 1 40768
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_48_387
timestamp 1698175906
transform 1 0 44688 0 1 40768
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_48_451
timestamp 1698175906
transform 1 0 51856 0 1 40768
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_48_457
timestamp 1698175906
transform 1 0 52528 0 1 40768
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_48_489
timestamp 1698175906
transform 1 0 56112 0 1 40768
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_48_505
timestamp 1698175906
transform 1 0 57904 0 1 40768
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_49_2
timestamp 1698175906
transform 1 0 1568 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_49_6
timestamp 1698175906
transform 1 0 2016 0 -1 42336
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_49_16
timestamp 1698175906
transform 1 0 3136 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_49_26
timestamp 1698175906
transform 1 0 4256 0 -1 42336
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_49_30
timestamp 1698175906
transform 1 0 4704 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_49_32
timestamp 1698175906
transform 1 0 4928 0 -1 42336
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_49_72
timestamp 1698175906
transform 1 0 9408 0 -1 42336
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_49_80
timestamp 1698175906
transform 1 0 10304 0 -1 42336
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_49_113
timestamp 1698175906
transform 1 0 14000 0 -1 42336
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_49_129
timestamp 1698175906
transform 1 0 15792 0 -1 42336
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_49_133
timestamp 1698175906
transform 1 0 16240 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_49_142
timestamp 1698175906
transform 1 0 17248 0 -1 42336
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_49_159
timestamp 1698175906
transform 1 0 19152 0 -1 42336
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_49_163
timestamp 1698175906
transform 1 0 19600 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_49_176
timestamp 1698175906
transform 1 0 21056 0 -1 42336
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_49_193
timestamp 1698175906
transform 1 0 22960 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_49_197
timestamp 1698175906
transform 1 0 23408 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_49_201
timestamp 1698175906
transform 1 0 23856 0 -1 42336
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_49_205
timestamp 1698175906
transform 1 0 24304 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_49_207
timestamp 1698175906
transform 1 0 24528 0 -1 42336
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_49_212
timestamp 1698175906
transform 1 0 25088 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_49_216
timestamp 1698175906
transform 1 0 25536 0 -1 42336
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_49_224
timestamp 1698175906
transform 1 0 26432 0 -1 42336
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_49_227
timestamp 1698175906
transform 1 0 26768 0 -1 42336
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_49_233
timestamp 1698175906
transform 1 0 27440 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_49_272
timestamp 1698175906
transform 1 0 31808 0 -1 42336
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_49_282
timestamp 1698175906
transform 1 0 32928 0 -1 42336
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_49_286
timestamp 1698175906
transform 1 0 33376 0 -1 42336
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_49_289
timestamp 1698175906
transform 1 0 33712 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_49_309
timestamp 1698175906
transform 1 0 35952 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_49_313
timestamp 1698175906
transform 1 0 36400 0 -1 42336
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_49_329
timestamp 1698175906
transform 1 0 38192 0 -1 42336
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_49_337
timestamp 1698175906
transform 1 0 39088 0 -1 42336
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_49_341
timestamp 1698175906
transform 1 0 39536 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_49_343
timestamp 1698175906
transform 1 0 39760 0 -1 42336
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_49_346
timestamp 1698175906
transform 1 0 40096 0 -1 42336
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_49_356
timestamp 1698175906
transform 1 0 41216 0 -1 42336
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_49_422
timestamp 1698175906
transform 1 0 48608 0 -1 42336
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_49_486
timestamp 1698175906
transform 1 0 55776 0 -1 42336
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_49_492
timestamp 1698175906
transform 1 0 56448 0 -1 42336
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_49_508
timestamp 1698175906
transform 1 0 58240 0 -1 42336
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_50_8
timestamp 1698175906
transform 1 0 2240 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_50_10
timestamp 1698175906
transform 1 0 2464 0 1 42336
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_50_16
timestamp 1698175906
transform 1 0 3136 0 1 42336
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_50_32
timestamp 1698175906
transform 1 0 4928 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_50_34
timestamp 1698175906
transform 1 0 5152 0 1 42336
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_50_37
timestamp 1698175906
transform 1 0 5488 0 1 42336
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_50_45
timestamp 1698175906
transform 1 0 6384 0 1 42336
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_50_49
timestamp 1698175906
transform 1 0 6832 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_50_102
timestamp 1698175906
transform 1 0 12768 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_50_104
timestamp 1698175906
transform 1 0 12992 0 1 42336
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_50_115
timestamp 1698175906
transform 1 0 14224 0 1 42336
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_50_131
timestamp 1698175906
transform 1 0 16016 0 1 42336
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_50_139
timestamp 1698175906
transform 1 0 16912 0 1 42336
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_50_143
timestamp 1698175906
transform 1 0 17360 0 1 42336
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_50_152
timestamp 1698175906
transform 1 0 18368 0 1 42336
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_50_168
timestamp 1698175906
transform 1 0 20160 0 1 42336
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_50_172
timestamp 1698175906
transform 1 0 20608 0 1 42336
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_50_185
timestamp 1698175906
transform 1 0 22064 0 1 42336
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_50_189
timestamp 1698175906
transform 1 0 22512 0 1 42336
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_50_192
timestamp 1698175906
transform 1 0 22848 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_50_196
timestamp 1698175906
transform 1 0 23296 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_50_239
timestamp 1698175906
transform 1 0 28112 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_50_243
timestamp 1698175906
transform 1 0 28560 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_50_247
timestamp 1698175906
transform 1 0 29008 0 1 42336
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_50_294
timestamp 1698175906
transform 1 0 34272 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_50_296
timestamp 1698175906
transform 1 0 34496 0 1 42336
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_50_299
timestamp 1698175906
transform 1 0 34832 0 1 42336
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_50_317
timestamp 1698175906
transform 1 0 36848 0 1 42336
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_50_325
timestamp 1698175906
transform 1 0 37744 0 1 42336
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_50_329
timestamp 1698175906
transform 1 0 38192 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_50_343
timestamp 1698175906
transform 1 0 39760 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_50_345
timestamp 1698175906
transform 1 0 39984 0 1 42336
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_50_383
timestamp 1698175906
transform 1 0 44240 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_50_387
timestamp 1698175906
transform 1 0 44688 0 1 42336
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_50_451
timestamp 1698175906
transform 1 0 51856 0 1 42336
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_50_457
timestamp 1698175906
transform 1 0 52528 0 1 42336
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_50_489
timestamp 1698175906
transform 1 0 56112 0 1 42336
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_50_505
timestamp 1698175906
transform 1 0 57904 0 1 42336
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_51_2
timestamp 1698175906
transform 1 0 1568 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_51_6
timestamp 1698175906
transform 1 0 2016 0 -1 43904
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_51_16
timestamp 1698175906
transform 1 0 3136 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_51_42
timestamp 1698175906
transform 1 0 6048 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_51_44
timestamp 1698175906
transform 1 0 6272 0 -1 43904
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_51_59
timestamp 1698175906
transform 1 0 7952 0 -1 43904
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_51_67
timestamp 1698175906
transform 1 0 8848 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_51_69
timestamp 1698175906
transform 1 0 9072 0 -1 43904
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_51_80
timestamp 1698175906
transform 1 0 10304 0 -1 43904
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_51_84
timestamp 1698175906
transform 1 0 10752 0 -1 43904
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_51_110
timestamp 1698175906
transform 1 0 13664 0 -1 43904
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_51_119
timestamp 1698175906
transform 1 0 14672 0 -1 43904
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_51_135
timestamp 1698175906
transform 1 0 16464 0 -1 43904
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_51_139
timestamp 1698175906
transform 1 0 16912 0 -1 43904
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_51_152
timestamp 1698175906
transform 1 0 18368 0 -1 43904
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_51_190
timestamp 1698175906
transform 1 0 22624 0 -1 43904
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_51_202
timestamp 1698175906
transform 1 0 23968 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_51_223
timestamp 1698175906
transform 1 0 26320 0 -1 43904
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_51_261
timestamp 1698175906
transform 1 0 30576 0 -1 43904
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_51_265
timestamp 1698175906
transform 1 0 31024 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_51_267
timestamp 1698175906
transform 1 0 31248 0 -1 43904
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_51_276
timestamp 1698175906
transform 1 0 32256 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_51_288
timestamp 1698175906
transform 1 0 33600 0 -1 43904
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_51_318
timestamp 1698175906
transform 1 0 36960 0 -1 43904
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_51_348
timestamp 1698175906
transform 1 0 40320 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_51_352
timestamp 1698175906
transform 1 0 40768 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_51_362
timestamp 1698175906
transform 1 0 41888 0 -1 43904
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_51_394
timestamp 1698175906
transform 1 0 45472 0 -1 43904
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_51_410
timestamp 1698175906
transform 1 0 47264 0 -1 43904
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_51_418
timestamp 1698175906
transform 1 0 48160 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_51_422
timestamp 1698175906
transform 1 0 48608 0 -1 43904
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_51_486
timestamp 1698175906
transform 1 0 55776 0 -1 43904
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_51_492
timestamp 1698175906
transform 1 0 56448 0 -1 43904
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_51_508
timestamp 1698175906
transform 1 0 58240 0 -1 43904
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_52_2
timestamp 1698175906
transform 1 0 1568 0 1 43904
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_52_34
timestamp 1698175906
transform 1 0 5152 0 1 43904
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_52_51
timestamp 1698175906
transform 1 0 7056 0 1 43904
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_52_67
timestamp 1698175906
transform 1 0 8848 0 1 43904
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_52_71
timestamp 1698175906
transform 1 0 9296 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_52_73
timestamp 1698175906
transform 1 0 9520 0 1 43904
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_52_98
timestamp 1698175906
transform 1 0 12320 0 1 43904
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_52_102
timestamp 1698175906
transform 1 0 12768 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_52_104
timestamp 1698175906
transform 1 0 12992 0 1 43904
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_52_107
timestamp 1698175906
transform 1 0 13328 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_52_109
timestamp 1698175906
transform 1 0 13552 0 1 43904
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_52_112
timestamp 1698175906
transform 1 0 13888 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_52_130
timestamp 1698175906
transform 1 0 15904 0 1 43904
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_52_187
timestamp 1698175906
transform 1 0 22288 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_52_189
timestamp 1698175906
transform 1 0 22512 0 1 43904
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_52_200
timestamp 1698175906
transform 1 0 23744 0 1 43904
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_52_231
timestamp 1698175906
transform 1 0 27216 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_52_257
timestamp 1698175906
transform 1 0 30128 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_52_259
timestamp 1698175906
transform 1 0 30352 0 1 43904
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_52_302
timestamp 1698175906
transform 1 0 35168 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_52_306
timestamp 1698175906
transform 1 0 35616 0 1 43904
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_52_314
timestamp 1698175906
transform 1 0 36512 0 1 43904
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_52_317
timestamp 1698175906
transform 1 0 36848 0 1 43904
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_52_325
timestamp 1698175906
transform 1 0 37744 0 1 43904
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_52_329
timestamp 1698175906
transform 1 0 38192 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_52_331
timestamp 1698175906
transform 1 0 38416 0 1 43904
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_52_342
timestamp 1698175906
transform 1 0 39648 0 1 43904
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_52_374
timestamp 1698175906
transform 1 0 43232 0 1 43904
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_52_382
timestamp 1698175906
transform 1 0 44128 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_52_384
timestamp 1698175906
transform 1 0 44352 0 1 43904
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_52_387
timestamp 1698175906
transform 1 0 44688 0 1 43904
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_52_451
timestamp 1698175906
transform 1 0 51856 0 1 43904
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_52_457
timestamp 1698175906
transform 1 0 52528 0 1 43904
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_52_489
timestamp 1698175906
transform 1 0 56112 0 1 43904
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_52_505
timestamp 1698175906
transform 1 0 57904 0 1 43904
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_53_2
timestamp 1698175906
transform 1 0 1568 0 -1 45472
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_53_6
timestamp 1698175906
transform 1 0 2016 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_53_8
timestamp 1698175906
transform 1 0 2240 0 -1 45472
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_53_19
timestamp 1698175906
transform 1 0 3472 0 -1 45472
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_53_28
timestamp 1698175906
transform 1 0 4480 0 -1 45472
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_53_64
timestamp 1698175906
transform 1 0 8512 0 -1 45472
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_53_68
timestamp 1698175906
transform 1 0 8960 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_53_72
timestamp 1698175906
transform 1 0 9408 0 -1 45472
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_53_99
timestamp 1698175906
transform 1 0 12432 0 -1 45472
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_53_107
timestamp 1698175906
transform 1 0 13328 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_53_109
timestamp 1698175906
transform 1 0 13552 0 -1 45472
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_53_118
timestamp 1698175906
transform 1 0 14560 0 -1 45472
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_53_134
timestamp 1698175906
transform 1 0 16352 0 -1 45472
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_53_138
timestamp 1698175906
transform 1 0 16800 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_53_142
timestamp 1698175906
transform 1 0 17248 0 -1 45472
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_53_150
timestamp 1698175906
transform 1 0 18144 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_53_152
timestamp 1698175906
transform 1 0 18368 0 -1 45472
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_53_199
timestamp 1698175906
transform 1 0 23632 0 -1 45472
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_53_203
timestamp 1698175906
transform 1 0 24080 0 -1 45472
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_53_206
timestamp 1698175906
transform 1 0 24416 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_53_212
timestamp 1698175906
transform 1 0 25088 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_53_214
timestamp 1698175906
transform 1 0 25312 0 -1 45472
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_53_257
timestamp 1698175906
transform 1 0 30128 0 -1 45472
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_53_273
timestamp 1698175906
transform 1 0 31920 0 -1 45472
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_53_277
timestamp 1698175906
transform 1 0 32368 0 -1 45472
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_53_282
timestamp 1698175906
transform 1 0 32928 0 -1 45472
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_53_339
timestamp 1698175906
transform 1 0 39312 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_53_341
timestamp 1698175906
transform 1 0 39536 0 -1 45472
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_53_352
timestamp 1698175906
transform 1 0 40768 0 -1 45472
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_53_356
timestamp 1698175906
transform 1 0 41216 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_53_387
timestamp 1698175906
transform 1 0 44688 0 -1 45472
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_53_419
timestamp 1698175906
transform 1 0 48272 0 -1 45472
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_53_422
timestamp 1698175906
transform 1 0 48608 0 -1 45472
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_53_486
timestamp 1698175906
transform 1 0 55776 0 -1 45472
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_53_492
timestamp 1698175906
transform 1 0 56448 0 -1 45472
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_53_508
timestamp 1698175906
transform 1 0 58240 0 -1 45472
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_54_8
timestamp 1698175906
transform 1 0 2240 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_54_12
timestamp 1698175906
transform 1 0 2688 0 1 45472
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_54_20
timestamp 1698175906
transform 1 0 3584 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_54_30
timestamp 1698175906
transform 1 0 4704 0 1 45472
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_54_34
timestamp 1698175906
transform 1 0 5152 0 1 45472
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_54_37
timestamp 1698175906
transform 1 0 5488 0 1 45472
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_54_67
timestamp 1698175906
transform 1 0 8848 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_54_69
timestamp 1698175906
transform 1 0 9072 0 1 45472
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_54_78
timestamp 1698175906
transform 1 0 10080 0 1 45472
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_54_107
timestamp 1698175906
transform 1 0 13328 0 1 45472
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_54_119
timestamp 1698175906
transform 1 0 14672 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_54_123
timestamp 1698175906
transform 1 0 15120 0 1 45472
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_54_127
timestamp 1698175906
transform 1 0 15568 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_54_129
timestamp 1698175906
transform 1 0 15792 0 1 45472
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_54_140
timestamp 1698175906
transform 1 0 17024 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_54_144
timestamp 1698175906
transform 1 0 17472 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_54_148
timestamp 1698175906
transform 1 0 17920 0 1 45472
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_54_156
timestamp 1698175906
transform 1 0 18816 0 1 45472
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_54_160
timestamp 1698175906
transform 1 0 19264 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_54_162
timestamp 1698175906
transform 1 0 19488 0 1 45472
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_54_169
timestamp 1698175906
transform 1 0 20272 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_54_173
timestamp 1698175906
transform 1 0 20720 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_54_191
timestamp 1698175906
transform 1 0 22736 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_54_287
timestamp 1698175906
transform 1 0 33488 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_54_291
timestamp 1698175906
transform 1 0 33936 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_54_301
timestamp 1698175906
transform 1 0 35056 0 1 45472
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_54_309
timestamp 1698175906
transform 1 0 35952 0 1 45472
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_54_313
timestamp 1698175906
transform 1 0 36400 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_54_317
timestamp 1698175906
transform 1 0 36848 0 1 45472
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_54_325
timestamp 1698175906
transform 1 0 37744 0 1 45472
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_54_329
timestamp 1698175906
transform 1 0 38192 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_54_335
timestamp 1698175906
transform 1 0 38864 0 1 45472
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_54_351
timestamp 1698175906
transform 1 0 40656 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_54_353
timestamp 1698175906
transform 1 0 40880 0 1 45472
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_54_364
timestamp 1698175906
transform 1 0 42112 0 1 45472
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_54_380
timestamp 1698175906
transform 1 0 43904 0 1 45472
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_54_384
timestamp 1698175906
transform 1 0 44352 0 1 45472
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_54_387
timestamp 1698175906
transform 1 0 44688 0 1 45472
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_54_451
timestamp 1698175906
transform 1 0 51856 0 1 45472
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_54_457
timestamp 1698175906
transform 1 0 52528 0 1 45472
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_54_489
timestamp 1698175906
transform 1 0 56112 0 1 45472
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_54_505
timestamp 1698175906
transform 1 0 57904 0 1 45472
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_55_8
timestamp 1698175906
transform 1 0 2240 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_55_12
timestamp 1698175906
transform 1 0 2688 0 -1 47040
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_55_26
timestamp 1698175906
transform 1 0 4256 0 -1 47040
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_55_72
timestamp 1698175906
transform 1 0 9408 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_55_126
timestamp 1698175906
transform 1 0 15456 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_55_130
timestamp 1698175906
transform 1 0 15904 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_55_134
timestamp 1698175906
transform 1 0 16352 0 -1 47040
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_55_138
timestamp 1698175906
transform 1 0 16800 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_55_142
timestamp 1698175906
transform 1 0 17248 0 -1 47040
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_55_158
timestamp 1698175906
transform 1 0 19040 0 -1 47040
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_55_162
timestamp 1698175906
transform 1 0 19488 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_55_164
timestamp 1698175906
transform 1 0 19712 0 -1 47040
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_55_171
timestamp 1698175906
transform 1 0 20496 0 -1 47040
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_55_187
timestamp 1698175906
transform 1 0 22288 0 -1 47040
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_55_193
timestamp 1698175906
transform 1 0 22960 0 -1 47040
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_55_201
timestamp 1698175906
transform 1 0 23856 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_55_203
timestamp 1698175906
transform 1 0 24080 0 -1 47040
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_55_206
timestamp 1698175906
transform 1 0 24416 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_55_262
timestamp 1698175906
transform 1 0 30688 0 -1 47040
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_55_290
timestamp 1698175906
transform 1 0 33824 0 -1 47040
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_55_294
timestamp 1698175906
transform 1 0 34272 0 -1 47040
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_55_324
timestamp 1698175906
transform 1 0 37632 0 -1 47040
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_55_332
timestamp 1698175906
transform 1 0 38528 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_55_342
timestamp 1698175906
transform 1 0 39648 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_55_346
timestamp 1698175906
transform 1 0 40096 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_55_360
timestamp 1698175906
transform 1 0 41664 0 -1 47040
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_55_392
timestamp 1698175906
transform 1 0 45248 0 -1 47040
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_55_408
timestamp 1698175906
transform 1 0 47040 0 -1 47040
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_55_416
timestamp 1698175906
transform 1 0 47936 0 -1 47040
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_55_422
timestamp 1698175906
transform 1 0 48608 0 -1 47040
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_55_486
timestamp 1698175906
transform 1 0 55776 0 -1 47040
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_55_492
timestamp 1698175906
transform 1 0 56448 0 -1 47040
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_55_508
timestamp 1698175906
transform 1 0 58240 0 -1 47040
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_56_2
timestamp 1698175906
transform 1 0 1568 0 1 47040
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_56_30
timestamp 1698175906
transform 1 0 4704 0 1 47040
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_56_34
timestamp 1698175906
transform 1 0 5152 0 1 47040
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_56_37
timestamp 1698175906
transform 1 0 5488 0 1 47040
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_56_41
timestamp 1698175906
transform 1 0 5936 0 1 47040
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_56_50
timestamp 1698175906
transform 1 0 6944 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_56_107
timestamp 1698175906
transform 1 0 13328 0 1 47040
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_56_132
timestamp 1698175906
transform 1 0 16128 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_56_136
timestamp 1698175906
transform 1 0 16576 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_56_145
timestamp 1698175906
transform 1 0 17584 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_56_147
timestamp 1698175906
transform 1 0 17808 0 1 47040
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_56_163
timestamp 1698175906
transform 1 0 19600 0 1 47040
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_56_171
timestamp 1698175906
transform 1 0 20496 0 1 47040
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_56_177
timestamp 1698175906
transform 1 0 21168 0 1 47040
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_56_193
timestamp 1698175906
transform 1 0 22960 0 1 47040
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_56_201
timestamp 1698175906
transform 1 0 23856 0 1 47040
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_56_205
timestamp 1698175906
transform 1 0 24304 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_56_207
timestamp 1698175906
transform 1 0 24528 0 1 47040
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_56_210
timestamp 1698175906
transform 1 0 24864 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_56_212
timestamp 1698175906
transform 1 0 25088 0 1 47040
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_56_279
timestamp 1698175906
transform 1 0 32592 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_56_305
timestamp 1698175906
transform 1 0 35504 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_56_309
timestamp 1698175906
transform 1 0 35952 0 1 47040
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_56_313
timestamp 1698175906
transform 1 0 36400 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_56_317
timestamp 1698175906
transform 1 0 36848 0 1 47040
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_56_333
timestamp 1698175906
transform 1 0 38640 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_56_372
timestamp 1698175906
transform 1 0 43008 0 1 47040
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_56_380
timestamp 1698175906
transform 1 0 43904 0 1 47040
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_56_384
timestamp 1698175906
transform 1 0 44352 0 1 47040
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_56_387
timestamp 1698175906
transform 1 0 44688 0 1 47040
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_56_451
timestamp 1698175906
transform 1 0 51856 0 1 47040
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_56_457
timestamp 1698175906
transform 1 0 52528 0 1 47040
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_56_489
timestamp 1698175906
transform 1 0 56112 0 1 47040
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_56_505
timestamp 1698175906
transform 1 0 57904 0 1 47040
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_57_2
timestamp 1698175906
transform 1 0 1568 0 -1 48608
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_57_26
timestamp 1698175906
transform 1 0 4256 0 -1 48608
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_57_34
timestamp 1698175906
transform 1 0 5152 0 -1 48608
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_57_38
timestamp 1698175906
transform 1 0 5600 0 -1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_57_40
timestamp 1698175906
transform 1 0 5824 0 -1 48608
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_57_54
timestamp 1698175906
transform 1 0 7392 0 -1 48608
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_57_72
timestamp 1698175906
transform 1 0 9408 0 -1 48608
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_57_97
timestamp 1698175906
transform 1 0 12208 0 -1 48608
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_57_105
timestamp 1698175906
transform 1 0 13104 0 -1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_57_107
timestamp 1698175906
transform 1 0 13328 0 -1 48608
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_57_118
timestamp 1698175906
transform 1 0 14560 0 -1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_57_130
timestamp 1698175906
transform 1 0 15904 0 -1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_57_134
timestamp 1698175906
transform 1 0 16352 0 -1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_57_138
timestamp 1698175906
transform 1 0 16800 0 -1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_57_142
timestamp 1698175906
transform 1 0 17248 0 -1 48608
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_57_170
timestamp 1698175906
transform 1 0 20384 0 -1 48608
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_57_178
timestamp 1698175906
transform 1 0 21280 0 -1 48608
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_57_185
timestamp 1698175906
transform 1 0 22064 0 -1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_57_187
timestamp 1698175906
transform 1 0 22288 0 -1 48608
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_57_205
timestamp 1698175906
transform 1 0 24304 0 -1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_57_209
timestamp 1698175906
transform 1 0 24752 0 -1 48608
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_57_212
timestamp 1698175906
transform 1 0 25088 0 -1 48608
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_57_220
timestamp 1698175906
transform 1 0 25984 0 -1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_57_222
timestamp 1698175906
transform 1 0 26208 0 -1 48608
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_57_273
timestamp 1698175906
transform 1 0 31920 0 -1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_57_277
timestamp 1698175906
transform 1 0 32368 0 -1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_57_279
timestamp 1698175906
transform 1 0 32592 0 -1 48608
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_57_282
timestamp 1698175906
transform 1 0 32928 0 -1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_57_284
timestamp 1698175906
transform 1 0 33152 0 -1 48608
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_57_343
timestamp 1698175906
transform 1 0 39760 0 -1 48608
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_57_347
timestamp 1698175906
transform 1 0 40208 0 -1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_57_349
timestamp 1698175906
transform 1 0 40432 0 -1 48608
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_57_352
timestamp 1698175906
transform 1 0 40768 0 -1 48608
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_57_416
timestamp 1698175906
transform 1 0 47936 0 -1 48608
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_57_422
timestamp 1698175906
transform 1 0 48608 0 -1 48608
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_57_486
timestamp 1698175906
transform 1 0 55776 0 -1 48608
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_57_492
timestamp 1698175906
transform 1 0 56448 0 -1 48608
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_57_508
timestamp 1698175906
transform 1 0 58240 0 -1 48608
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_58_8
timestamp 1698175906
transform 1 0 2240 0 1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_58_12
timestamp 1698175906
transform 1 0 2688 0 1 48608
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_58_28
timestamp 1698175906
transform 1 0 4480 0 1 48608
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_58_32
timestamp 1698175906
transform 1 0 4928 0 1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_58_34
timestamp 1698175906
transform 1 0 5152 0 1 48608
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_58_37
timestamp 1698175906
transform 1 0 5488 0 1 48608
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_58_53
timestamp 1698175906
transform 1 0 7280 0 1 48608
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_58_69
timestamp 1698175906
transform 1 0 9072 0 1 48608
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_58_81
timestamp 1698175906
transform 1 0 10416 0 1 48608
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_58_85
timestamp 1698175906
transform 1 0 10864 0 1 48608
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_58_92
timestamp 1698175906
transform 1 0 11648 0 1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_58_96
timestamp 1698175906
transform 1 0 12096 0 1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_58_98
timestamp 1698175906
transform 1 0 12320 0 1 48608
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_58_101
timestamp 1698175906
transform 1 0 12656 0 1 48608
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_58_107
timestamp 1698175906
transform 1 0 13328 0 1 48608
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_58_115
timestamp 1698175906
transform 1 0 14224 0 1 48608
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_58_118
timestamp 1698175906
transform 1 0 14560 0 1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_58_137
timestamp 1698175906
transform 1 0 16688 0 1 48608
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_58_145
timestamp 1698175906
transform 1 0 17584 0 1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_58_147
timestamp 1698175906
transform 1 0 17808 0 1 48608
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_58_160
timestamp 1698175906
transform 1 0 19264 0 1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_58_164
timestamp 1698175906
transform 1 0 19712 0 1 48608
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_58_173
timestamp 1698175906
transform 1 0 20720 0 1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_58_177
timestamp 1698175906
transform 1 0 21168 0 1 48608
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_58_196
timestamp 1698175906
transform 1 0 23296 0 1 48608
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_58_204
timestamp 1698175906
transform 1 0 24192 0 1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_58_242
timestamp 1698175906
transform 1 0 28448 0 1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_58_244
timestamp 1698175906
transform 1 0 28672 0 1 48608
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_58_247
timestamp 1698175906
transform 1 0 29008 0 1 48608
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_58_280
timestamp 1698175906
transform 1 0 32704 0 1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_58_284
timestamp 1698175906
transform 1 0 33152 0 1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_58_317
timestamp 1698175906
transform 1 0 36848 0 1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_58_321
timestamp 1698175906
transform 1 0 37296 0 1 48608
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_58_329
timestamp 1698175906
transform 1 0 38192 0 1 48608
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_58_333
timestamp 1698175906
transform 1 0 38640 0 1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_58_337
timestamp 1698175906
transform 1 0 39088 0 1 48608
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_58_369
timestamp 1698175906
transform 1 0 42672 0 1 48608
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_58_387
timestamp 1698175906
transform 1 0 44688 0 1 48608
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_58_451
timestamp 1698175906
transform 1 0 51856 0 1 48608
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_58_457
timestamp 1698175906
transform 1 0 52528 0 1 48608
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_58_489
timestamp 1698175906
transform 1 0 56112 0 1 48608
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_58_505
timestamp 1698175906
transform 1 0 57904 0 1 48608
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_59_31
timestamp 1698175906
transform 1 0 4816 0 -1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_59_35
timestamp 1698175906
transform 1 0 5264 0 -1 50176
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_59_39
timestamp 1698175906
transform 1 0 5712 0 -1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_59_41
timestamp 1698175906
transform 1 0 5936 0 -1 50176
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_59_72
timestamp 1698175906
transform 1 0 9408 0 -1 50176
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_59_84
timestamp 1698175906
transform 1 0 10752 0 -1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_59_86
timestamp 1698175906
transform 1 0 10976 0 -1 50176
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_59_99
timestamp 1698175906
transform 1 0 12432 0 -1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_59_107
timestamp 1698175906
transform 1 0 13328 0 -1 50176
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_59_139
timestamp 1698175906
transform 1 0 16912 0 -1 50176
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_59_192
timestamp 1698175906
transform 1 0 22848 0 -1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_59_196
timestamp 1698175906
transform 1 0 23296 0 -1 50176
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_59_200
timestamp 1698175906
transform 1 0 23744 0 -1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_59_202
timestamp 1698175906
transform 1 0 23968 0 -1 50176
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_59_205
timestamp 1698175906
transform 1 0 24304 0 -1 50176
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_59_209
timestamp 1698175906
transform 1 0 24752 0 -1 50176
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_59_216
timestamp 1698175906
transform 1 0 25536 0 -1 50176
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_59_232
timestamp 1698175906
transform 1 0 27328 0 -1 50176
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_59_237
timestamp 1698175906
transform 1 0 27888 0 -1 50176
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_59_245
timestamp 1698175906
transform 1 0 28784 0 -1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_59_247
timestamp 1698175906
transform 1 0 29008 0 -1 50176
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_59_277
timestamp 1698175906
transform 1 0 32368 0 -1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_59_279
timestamp 1698175906
transform 1 0 32592 0 -1 50176
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_59_290
timestamp 1698175906
transform 1 0 33824 0 -1 50176
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_59_302
timestamp 1698175906
transform 1 0 35168 0 -1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_59_306
timestamp 1698175906
transform 1 0 35616 0 -1 50176
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_59_338
timestamp 1698175906
transform 1 0 39200 0 -1 50176
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_59_346
timestamp 1698175906
transform 1 0 40096 0 -1 50176
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_59_352
timestamp 1698175906
transform 1 0 40768 0 -1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_59_356
timestamp 1698175906
transform 1 0 41216 0 -1 50176
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_59_422
timestamp 1698175906
transform 1 0 48608 0 -1 50176
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_59_486
timestamp 1698175906
transform 1 0 55776 0 -1 50176
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_59_492
timestamp 1698175906
transform 1 0 56448 0 -1 50176
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_59_508
timestamp 1698175906
transform 1 0 58240 0 -1 50176
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_60_31
timestamp 1698175906
transform 1 0 4816 0 1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_60_37
timestamp 1698175906
transform 1 0 5488 0 1 50176
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_60_45
timestamp 1698175906
transform 1 0 6384 0 1 50176
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_60_49
timestamp 1698175906
transform 1 0 6832 0 1 50176
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_60_58
timestamp 1698175906
transform 1 0 7840 0 1 50176
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_60_90
timestamp 1698175906
transform 1 0 11424 0 1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_60_92
timestamp 1698175906
transform 1 0 11648 0 1 50176
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_60_95
timestamp 1698175906
transform 1 0 11984 0 1 50176
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_60_101
timestamp 1698175906
transform 1 0 12656 0 1 50176
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_60_107
timestamp 1698175906
transform 1 0 13328 0 1 50176
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_60_123
timestamp 1698175906
transform 1 0 15120 0 1 50176
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_60_127
timestamp 1698175906
transform 1 0 15568 0 1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_60_133
timestamp 1698175906
transform 1 0 16240 0 1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_60_137
timestamp 1698175906
transform 1 0 16688 0 1 50176
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_60_145
timestamp 1698175906
transform 1 0 17584 0 1 50176
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_60_154
timestamp 1698175906
transform 1 0 18592 0 1 50176
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_60_170
timestamp 1698175906
transform 1 0 20384 0 1 50176
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_60_174
timestamp 1698175906
transform 1 0 20832 0 1 50176
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_60_177
timestamp 1698175906
transform 1 0 21168 0 1 50176
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_60_181
timestamp 1698175906
transform 1 0 21616 0 1 50176
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_60_190
timestamp 1698175906
transform 1 0 22624 0 1 50176
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_60_194
timestamp 1698175906
transform 1 0 23072 0 1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_60_196
timestamp 1698175906
transform 1 0 23296 0 1 50176
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_60_211
timestamp 1698175906
transform 1 0 24976 0 1 50176
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_60_219
timestamp 1698175906
transform 1 0 25872 0 1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_60_221
timestamp 1698175906
transform 1 0 26096 0 1 50176
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_60_230
timestamp 1698175906
transform 1 0 27104 0 1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_60_234
timestamp 1698175906
transform 1 0 27552 0 1 50176
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_60_242
timestamp 1698175906
transform 1 0 28448 0 1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_60_244
timestamp 1698175906
transform 1 0 28672 0 1 50176
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_60_247
timestamp 1698175906
transform 1 0 29008 0 1 50176
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_60_255
timestamp 1698175906
transform 1 0 29904 0 1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_60_257
timestamp 1698175906
transform 1 0 30128 0 1 50176
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_60_264
timestamp 1698175906
transform 1 0 30912 0 1 50176
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_60_272
timestamp 1698175906
transform 1 0 31808 0 1 50176
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_60_276
timestamp 1698175906
transform 1 0 32256 0 1 50176
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_60_279
timestamp 1698175906
transform 1 0 32592 0 1 50176
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_60_295
timestamp 1698175906
transform 1 0 34384 0 1 50176
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_60_304
timestamp 1698175906
transform 1 0 35392 0 1 50176
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_60_312
timestamp 1698175906
transform 1 0 36288 0 1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_60_314
timestamp 1698175906
transform 1 0 36512 0 1 50176
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_60_317
timestamp 1698175906
transform 1 0 36848 0 1 50176
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_60_347
timestamp 1698175906
transform 1 0 40208 0 1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_60_351
timestamp 1698175906
transform 1 0 40656 0 1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_60_384
timestamp 1698175906
transform 1 0 44352 0 1 50176
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_60_387
timestamp 1698175906
transform 1 0 44688 0 1 50176
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_60_451
timestamp 1698175906
transform 1 0 51856 0 1 50176
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_60_457
timestamp 1698175906
transform 1 0 52528 0 1 50176
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_60_489
timestamp 1698175906
transform 1 0 56112 0 1 50176
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_60_505
timestamp 1698175906
transform 1 0 57904 0 1 50176
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_61_8
timestamp 1698175906
transform 1 0 2240 0 -1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_61_12
timestamp 1698175906
transform 1 0 2688 0 -1 51744
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_61_20
timestamp 1698175906
transform 1 0 3584 0 -1 51744
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_61_24
timestamp 1698175906
transform 1 0 4032 0 -1 51744
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_61_54
timestamp 1698175906
transform 1 0 7392 0 -1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_61_58
timestamp 1698175906
transform 1 0 7840 0 -1 51744
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_61_66
timestamp 1698175906
transform 1 0 8736 0 -1 51744
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_61_72
timestamp 1698175906
transform 1 0 9408 0 -1 51744
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_61_80
timestamp 1698175906
transform 1 0 10304 0 -1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_61_92
timestamp 1698175906
transform 1 0 11648 0 -1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_61_96
timestamp 1698175906
transform 1 0 12096 0 -1 51744
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_61_133
timestamp 1698175906
transform 1 0 16240 0 -1 51744
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_61_148
timestamp 1698175906
transform 1 0 17920 0 -1 51744
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_61_157
timestamp 1698175906
transform 1 0 18928 0 -1 51744
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_61_173
timestamp 1698175906
transform 1 0 20720 0 -1 51744
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_61_203
timestamp 1698175906
transform 1 0 24080 0 -1 51744
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_61_207
timestamp 1698175906
transform 1 0 24528 0 -1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_61_209
timestamp 1698175906
transform 1 0 24752 0 -1 51744
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_61_212
timestamp 1698175906
transform 1 0 25088 0 -1 51744
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_61_242
timestamp 1698175906
transform 1 0 28448 0 -1 51744
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_61_274
timestamp 1698175906
transform 1 0 32032 0 -1 51744
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_61_278
timestamp 1698175906
transform 1 0 32480 0 -1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_61_282
timestamp 1698175906
transform 1 0 32928 0 -1 51744
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_61_314
timestamp 1698175906
transform 1 0 36512 0 -1 51744
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_61_330
timestamp 1698175906
transform 1 0 38304 0 -1 51744
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_61_349
timestamp 1698175906
transform 1 0 40432 0 -1 51744
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_61_352
timestamp 1698175906
transform 1 0 40768 0 -1 51744
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_61_369
timestamp 1698175906
transform 1 0 42672 0 -1 51744
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_61_401
timestamp 1698175906
transform 1 0 46256 0 -1 51744
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_61_417
timestamp 1698175906
transform 1 0 48048 0 -1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_61_419
timestamp 1698175906
transform 1 0 48272 0 -1 51744
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_61_422
timestamp 1698175906
transform 1 0 48608 0 -1 51744
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_61_486
timestamp 1698175906
transform 1 0 55776 0 -1 51744
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_61_492
timestamp 1698175906
transform 1 0 56448 0 -1 51744
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_61_508
timestamp 1698175906
transform 1 0 58240 0 -1 51744
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_62_2
timestamp 1698175906
transform 1 0 1568 0 1 51744
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_62_34
timestamp 1698175906
transform 1 0 5152 0 1 51744
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_62_37
timestamp 1698175906
transform 1 0 5488 0 1 51744
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_62_53
timestamp 1698175906
transform 1 0 7280 0 1 51744
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_62_61
timestamp 1698175906
transform 1 0 8176 0 1 51744
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_62_65
timestamp 1698175906
transform 1 0 8624 0 1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_62_67
timestamp 1698175906
transform 1 0 8848 0 1 51744
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_62_70
timestamp 1698175906
transform 1 0 9184 0 1 51744
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_62_74
timestamp 1698175906
transform 1 0 9632 0 1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_62_96
timestamp 1698175906
transform 1 0 12096 0 1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_62_100
timestamp 1698175906
transform 1 0 12544 0 1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_62_104
timestamp 1698175906
transform 1 0 12992 0 1 51744
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_62_107
timestamp 1698175906
transform 1 0 13328 0 1 51744
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_62_115
timestamp 1698175906
transform 1 0 14224 0 1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_62_125
timestamp 1698175906
transform 1 0 15344 0 1 51744
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_62_134
timestamp 1698175906
transform 1 0 16352 0 1 51744
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_62_142
timestamp 1698175906
transform 1 0 17248 0 1 51744
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_62_177
timestamp 1698175906
transform 1 0 21168 0 1 51744
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_62_181
timestamp 1698175906
transform 1 0 21616 0 1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_62_233
timestamp 1698175906
transform 1 0 27440 0 1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_62_237
timestamp 1698175906
transform 1 0 27888 0 1 51744
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_62_247
timestamp 1698175906
transform 1 0 29008 0 1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_62_278
timestamp 1698175906
transform 1 0 32480 0 1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_62_280
timestamp 1698175906
transform 1 0 32704 0 1 51744
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_62_283
timestamp 1698175906
transform 1 0 33040 0 1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_62_314
timestamp 1698175906
transform 1 0 36512 0 1 51744
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_62_317
timestamp 1698175906
transform 1 0 36848 0 1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_62_321
timestamp 1698175906
transform 1 0 37296 0 1 51744
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_62_379
timestamp 1698175906
transform 1 0 43792 0 1 51744
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_62_383
timestamp 1698175906
transform 1 0 44240 0 1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_62_387
timestamp 1698175906
transform 1 0 44688 0 1 51744
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_62_451
timestamp 1698175906
transform 1 0 51856 0 1 51744
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_62_457
timestamp 1698175906
transform 1 0 52528 0 1 51744
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_62_489
timestamp 1698175906
transform 1 0 56112 0 1 51744
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_62_505
timestamp 1698175906
transform 1 0 57904 0 1 51744
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_63_8
timestamp 1698175906
transform 1 0 2240 0 -1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_63_12
timestamp 1698175906
transform 1 0 2688 0 -1 53312
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_63_28
timestamp 1698175906
transform 1 0 4480 0 -1 53312
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_63_36
timestamp 1698175906
transform 1 0 5376 0 -1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_63_38
timestamp 1698175906
transform 1 0 5600 0 -1 53312
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_63_68
timestamp 1698175906
transform 1 0 8960 0 -1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_63_72
timestamp 1698175906
transform 1 0 9408 0 -1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_63_74
timestamp 1698175906
transform 1 0 9632 0 -1 53312
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_63_91
timestamp 1698175906
transform 1 0 11536 0 -1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_63_93
timestamp 1698175906
transform 1 0 11760 0 -1 53312
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_63_100
timestamp 1698175906
transform 1 0 12544 0 -1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_63_104
timestamp 1698175906
transform 1 0 12992 0 -1 53312
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_63_120
timestamp 1698175906
transform 1 0 14784 0 -1 53312
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_63_124
timestamp 1698175906
transform 1 0 15232 0 -1 53312
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_63_127
timestamp 1698175906
transform 1 0 15568 0 -1 53312
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_63_135
timestamp 1698175906
transform 1 0 16464 0 -1 53312
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_63_139
timestamp 1698175906
transform 1 0 16912 0 -1 53312
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_63_142
timestamp 1698175906
transform 1 0 17248 0 -1 53312
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_63_146
timestamp 1698175906
transform 1 0 17696 0 -1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_63_156
timestamp 1698175906
transform 1 0 18816 0 -1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_63_160
timestamp 1698175906
transform 1 0 19264 0 -1 53312
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_63_176
timestamp 1698175906
transform 1 0 21056 0 -1 53312
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_63_184
timestamp 1698175906
transform 1 0 21952 0 -1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_63_186
timestamp 1698175906
transform 1 0 22176 0 -1 53312
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_63_195
timestamp 1698175906
transform 1 0 23184 0 -1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_63_199
timestamp 1698175906
transform 1 0 23632 0 -1 53312
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_63_207
timestamp 1698175906
transform 1 0 24528 0 -1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_63_209
timestamp 1698175906
transform 1 0 24752 0 -1 53312
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_63_212
timestamp 1698175906
transform 1 0 25088 0 -1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_63_214
timestamp 1698175906
transform 1 0 25312 0 -1 53312
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_63_223
timestamp 1698175906
transform 1 0 26320 0 -1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_63_231
timestamp 1698175906
transform 1 0 27216 0 -1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_63_235
timestamp 1698175906
transform 1 0 27664 0 -1 53312
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_63_243
timestamp 1698175906
transform 1 0 28560 0 -1 53312
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_63_247
timestamp 1698175906
transform 1 0 29008 0 -1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_63_265
timestamp 1698175906
transform 1 0 31024 0 -1 53312
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_63_269
timestamp 1698175906
transform 1 0 31472 0 -1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_63_271
timestamp 1698175906
transform 1 0 31696 0 -1 53312
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_63_278
timestamp 1698175906
transform 1 0 32480 0 -1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_63_282
timestamp 1698175906
transform 1 0 32928 0 -1 53312
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_63_293
timestamp 1698175906
transform 1 0 34160 0 -1 53312
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_63_309
timestamp 1698175906
transform 1 0 35952 0 -1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_63_311
timestamp 1698175906
transform 1 0 36176 0 -1 53312
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_63_329
timestamp 1698175906
transform 1 0 38192 0 -1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_63_333
timestamp 1698175906
transform 1 0 38640 0 -1 53312
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_63_349
timestamp 1698175906
transform 1 0 40432 0 -1 53312
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_63_352
timestamp 1698175906
transform 1 0 40768 0 -1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_63_356
timestamp 1698175906
transform 1 0 41216 0 -1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_63_358
timestamp 1698175906
transform 1 0 41440 0 -1 53312
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_63_390
timestamp 1698175906
transform 1 0 45024 0 -1 53312
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_63_406
timestamp 1698175906
transform 1 0 46816 0 -1 53312
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_63_414
timestamp 1698175906
transform 1 0 47712 0 -1 53312
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_63_418
timestamp 1698175906
transform 1 0 48160 0 -1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_63_422
timestamp 1698175906
transform 1 0 48608 0 -1 53312
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_63_486
timestamp 1698175906
transform 1 0 55776 0 -1 53312
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_63_492
timestamp 1698175906
transform 1 0 56448 0 -1 53312
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_63_508
timestamp 1698175906
transform 1 0 58240 0 -1 53312
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_64_2
timestamp 1698175906
transform 1 0 1568 0 1 53312
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_64_34
timestamp 1698175906
transform 1 0 5152 0 1 53312
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_64_37
timestamp 1698175906
transform 1 0 5488 0 1 53312
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_64_69
timestamp 1698175906
transform 1 0 9072 0 1 53312
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_64_77
timestamp 1698175906
transform 1 0 9968 0 1 53312
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_64_83
timestamp 1698175906
transform 1 0 10640 0 1 53312
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_64_93
timestamp 1698175906
transform 1 0 11760 0 1 53312
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_64_101
timestamp 1698175906
transform 1 0 12656 0 1 53312
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_64_107
timestamp 1698175906
transform 1 0 13328 0 1 53312
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_64_123
timestamp 1698175906
transform 1 0 15120 0 1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_64_125
timestamp 1698175906
transform 1 0 15344 0 1 53312
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_64_128
timestamp 1698175906
transform 1 0 15680 0 1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_64_130
timestamp 1698175906
transform 1 0 15904 0 1 53312
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_64_139
timestamp 1698175906
transform 1 0 16912 0 1 53312
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_64_147
timestamp 1698175906
transform 1 0 17808 0 1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_64_149
timestamp 1698175906
transform 1 0 18032 0 1 53312
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_64_152
timestamp 1698175906
transform 1 0 18368 0 1 53312
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_64_168
timestamp 1698175906
transform 1 0 20160 0 1 53312
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_64_172
timestamp 1698175906
transform 1 0 20608 0 1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_64_174
timestamp 1698175906
transform 1 0 20832 0 1 53312
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_64_177
timestamp 1698175906
transform 1 0 21168 0 1 53312
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_64_181
timestamp 1698175906
transform 1 0 21616 0 1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_64_183
timestamp 1698175906
transform 1 0 21840 0 1 53312
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_64_194
timestamp 1698175906
transform 1 0 23072 0 1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_64_196
timestamp 1698175906
transform 1 0 23296 0 1 53312
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_64_205
timestamp 1698175906
transform 1 0 24304 0 1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_64_215
timestamp 1698175906
transform 1 0 25424 0 1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_64_219
timestamp 1698175906
transform 1 0 25872 0 1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_64_229
timestamp 1698175906
transform 1 0 26992 0 1 53312
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_64_247
timestamp 1698175906
transform 1 0 29008 0 1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_64_251
timestamp 1698175906
transform 1 0 29456 0 1 53312
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_64_267
timestamp 1698175906
transform 1 0 31248 0 1 53312
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_64_275
timestamp 1698175906
transform 1 0 32144 0 1 53312
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_64_287
timestamp 1698175906
transform 1 0 33488 0 1 53312
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_64_303
timestamp 1698175906
transform 1 0 35280 0 1 53312
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_64_311
timestamp 1698175906
transform 1 0 36176 0 1 53312
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_64_317
timestamp 1698175906
transform 1 0 36848 0 1 53312
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_64_339
timestamp 1698175906
transform 1 0 39312 0 1 53312
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_64_347
timestamp 1698175906
transform 1 0 40208 0 1 53312
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_64_351
timestamp 1698175906
transform 1 0 40656 0 1 53312
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_64_358
timestamp 1698175906
transform 1 0 41440 0 1 53312
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_64_362
timestamp 1698175906
transform 1 0 41888 0 1 53312
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_64_369
timestamp 1698175906
transform 1 0 42672 0 1 53312
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_64_387
timestamp 1698175906
transform 1 0 44688 0 1 53312
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_64_451
timestamp 1698175906
transform 1 0 51856 0 1 53312
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_64_457
timestamp 1698175906
transform 1 0 52528 0 1 53312
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_64_489
timestamp 1698175906
transform 1 0 56112 0 1 53312
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_64_505
timestamp 1698175906
transform 1 0 57904 0 1 53312
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_65_8
timestamp 1698175906
transform 1 0 2240 0 -1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_65_12
timestamp 1698175906
transform 1 0 2688 0 -1 54880
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_65_44
timestamp 1698175906
transform 1 0 6272 0 -1 54880
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_65_60
timestamp 1698175906
transform 1 0 8064 0 -1 54880
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_65_68
timestamp 1698175906
transform 1 0 8960 0 -1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_65_72
timestamp 1698175906
transform 1 0 9408 0 -1 54880
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_65_88
timestamp 1698175906
transform 1 0 11200 0 -1 54880
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_65_96
timestamp 1698175906
transform 1 0 12096 0 -1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_65_113
timestamp 1698175906
transform 1 0 14000 0 -1 54880
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_65_117
timestamp 1698175906
transform 1 0 14448 0 -1 54880
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_65_126
timestamp 1698175906
transform 1 0 15456 0 -1 54880
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_65_135
timestamp 1698175906
transform 1 0 16464 0 -1 54880
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_65_139
timestamp 1698175906
transform 1 0 16912 0 -1 54880
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_65_158
timestamp 1698175906
transform 1 0 19040 0 -1 54880
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_65_203
timestamp 1698175906
transform 1 0 24080 0 -1 54880
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_65_207
timestamp 1698175906
transform 1 0 24528 0 -1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_65_209
timestamp 1698175906
transform 1 0 24752 0 -1 54880
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_65_241
timestamp 1698175906
transform 1 0 28336 0 -1 54880
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_65_263
timestamp 1698175906
transform 1 0 30800 0 -1 54880
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_65_267
timestamp 1698175906
transform 1 0 31248 0 -1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_65_269
timestamp 1698175906
transform 1 0 31472 0 -1 54880
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_65_276
timestamp 1698175906
transform 1 0 32256 0 -1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_65_282
timestamp 1698175906
transform 1 0 32928 0 -1 54880
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_65_293
timestamp 1698175906
transform 1 0 34160 0 -1 54880
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_65_300
timestamp 1698175906
transform 1 0 34944 0 -1 54880
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_65_308
timestamp 1698175906
transform 1 0 35840 0 -1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_65_310
timestamp 1698175906
transform 1 0 36064 0 -1 54880
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_65_317
timestamp 1698175906
transform 1 0 36848 0 -1 54880
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_65_325
timestamp 1698175906
transform 1 0 37744 0 -1 54880
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_65_337
timestamp 1698175906
transform 1 0 39088 0 -1 54880
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_65_345
timestamp 1698175906
transform 1 0 39984 0 -1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_65_347
timestamp 1698175906
transform 1 0 40208 0 -1 54880
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_65_362
timestamp 1698175906
transform 1 0 41888 0 -1 54880
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_65_394
timestamp 1698175906
transform 1 0 45472 0 -1 54880
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_65_410
timestamp 1698175906
transform 1 0 47264 0 -1 54880
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_65_418
timestamp 1698175906
transform 1 0 48160 0 -1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_65_422
timestamp 1698175906
transform 1 0 48608 0 -1 54880
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_65_454
timestamp 1698175906
transform 1 0 52192 0 -1 54880
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_65_470
timestamp 1698175906
transform 1 0 53984 0 -1 54880
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_65_478
timestamp 1698175906
transform 1 0 54880 0 -1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_65_480
timestamp 1698175906
transform 1 0 55104 0 -1 54880
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_65_483
timestamp 1698175906
transform 1 0 55440 0 -1 54880
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_65_487
timestamp 1698175906
transform 1 0 55888 0 -1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_65_489
timestamp 1698175906
transform 1 0 56112 0 -1 54880
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_65_492
timestamp 1698175906
transform 1 0 56448 0 -1 54880
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_65_508
timestamp 1698175906
transform 1 0 58240 0 -1 54880
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_66_2
timestamp 1698175906
transform 1 0 1568 0 1 54880
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_66_8
timestamp 1698175906
transform 1 0 2240 0 1 54880
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_66_24
timestamp 1698175906
transform 1 0 4032 0 1 54880
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_66_32
timestamp 1698175906
transform 1 0 4928 0 1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_66_34
timestamp 1698175906
transform 1 0 5152 0 1 54880
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_66_37
timestamp 1698175906
transform 1 0 5488 0 1 54880
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_66_69
timestamp 1698175906
transform 1 0 9072 0 1 54880
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_66_85
timestamp 1698175906
transform 1 0 10864 0 1 54880
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_66_89
timestamp 1698175906
transform 1 0 11312 0 1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_66_91
timestamp 1698175906
transform 1 0 11536 0 1 54880
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_66_96
timestamp 1698175906
transform 1 0 12096 0 1 54880
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_66_104
timestamp 1698175906
transform 1 0 12992 0 1 54880
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_66_136
timestamp 1698175906
transform 1 0 16576 0 1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_66_140
timestamp 1698175906
transform 1 0 17024 0 1 54880
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_66_173
timestamp 1698175906
transform 1 0 20720 0 1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_66_177
timestamp 1698175906
transform 1 0 21168 0 1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_66_181
timestamp 1698175906
transform 1 0 21616 0 1 54880
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_66_189
timestamp 1698175906
transform 1 0 22512 0 1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_66_195
timestamp 1698175906
transform 1 0 23184 0 1 54880
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_66_211
timestamp 1698175906
transform 1 0 24976 0 1 54880
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_66_216
timestamp 1698175906
transform 1 0 25536 0 1 54880
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_66_232
timestamp 1698175906
transform 1 0 27328 0 1 54880
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_66_237
timestamp 1698175906
transform 1 0 27888 0 1 54880
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_66_282
timestamp 1698175906
transform 1 0 32928 0 1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_66_323
timestamp 1698175906
transform 1 0 37520 0 1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_66_327
timestamp 1698175906
transform 1 0 37968 0 1 54880
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_66_340
timestamp 1698175906
transform 1 0 39424 0 1 54880
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_66_375
timestamp 1698175906
transform 1 0 43344 0 1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_66_379
timestamp 1698175906
transform 1 0 43792 0 1 54880
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_66_383
timestamp 1698175906
transform 1 0 44240 0 1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_66_387
timestamp 1698175906
transform 1 0 44688 0 1 54880
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_66_391
timestamp 1698175906
transform 1 0 45136 0 1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_66_421
timestamp 1698175906
transform 1 0 48496 0 1 54880
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_66_437
timestamp 1698175906
transform 1 0 50288 0 1 54880
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_66_441
timestamp 1698175906
transform 1 0 50736 0 1 54880
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_66_444
timestamp 1698175906
transform 1 0 51072 0 1 54880
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_66_452
timestamp 1698175906
transform 1 0 51968 0 1 54880
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_67_14
timestamp 1698175906
transform 1 0 2912 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_67_18
timestamp 1698175906
transform 1 0 3360 0 -1 56448
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_67_26
timestamp 1698175906
transform 1 0 4256 0 -1 56448
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_67_30
timestamp 1698175906
transform 1 0 4704 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_67_42
timestamp 1698175906
transform 1 0 6048 0 -1 56448
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_67_50
timestamp 1698175906
transform 1 0 6944 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_67_52
timestamp 1698175906
transform 1 0 7168 0 -1 56448
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_67_61
timestamp 1698175906
transform 1 0 8176 0 -1 56448
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_67_65
timestamp 1698175906
transform 1 0 8624 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_67_67
timestamp 1698175906
transform 1 0 8848 0 -1 56448
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_67_70
timestamp 1698175906
transform 1 0 9184 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_67_72
timestamp 1698175906
transform 1 0 9408 0 -1 56448
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_67_81
timestamp 1698175906
transform 1 0 10416 0 -1 56448
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_67_89
timestamp 1698175906
transform 1 0 11312 0 -1 56448
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_67_101
timestamp 1698175906
transform 1 0 12656 0 -1 56448
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_67_104
timestamp 1698175906
transform 1 0 12992 0 -1 56448
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_67_112
timestamp 1698175906
transform 1 0 13888 0 -1 56448
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_67_121
timestamp 1698175906
transform 1 0 14896 0 -1 56448
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_67_129
timestamp 1698175906
transform 1 0 15792 0 -1 56448
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_67_133
timestamp 1698175906
transform 1 0 16240 0 -1 56448
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_67_144
timestamp 1698175906
transform 1 0 17472 0 -1 56448
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_67_152
timestamp 1698175906
transform 1 0 18368 0 -1 56448
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_67_161
timestamp 1698175906
transform 1 0 19376 0 -1 56448
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_67_165
timestamp 1698175906
transform 1 0 19824 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_67_167
timestamp 1698175906
transform 1 0 20048 0 -1 56448
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_67_172
timestamp 1698175906
transform 1 0 20608 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_67_174
timestamp 1698175906
transform 1 0 20832 0 -1 56448
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_67_181
timestamp 1698175906
transform 1 0 21616 0 -1 56448
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_67_189
timestamp 1698175906
transform 1 0 22512 0 -1 56448
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_67_201
timestamp 1698175906
transform 1 0 23856 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_67_203
timestamp 1698175906
transform 1 0 24080 0 -1 56448
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_67_206
timestamp 1698175906
transform 1 0 24416 0 -1 56448
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_67_210
timestamp 1698175906
transform 1 0 24864 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_67_212
timestamp 1698175906
transform 1 0 25088 0 -1 56448
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_67_221
timestamp 1698175906
transform 1 0 26096 0 -1 56448
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_67_229
timestamp 1698175906
transform 1 0 26992 0 -1 56448
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_67_233
timestamp 1698175906
transform 1 0 27440 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_67_235
timestamp 1698175906
transform 1 0 27664 0 -1 56448
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_67_246
timestamp 1698175906
transform 1 0 28896 0 -1 56448
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_67_250
timestamp 1698175906
transform 1 0 29344 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_67_252
timestamp 1698175906
transform 1 0 29568 0 -1 56448
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_67_261
timestamp 1698175906
transform 1 0 30576 0 -1 56448
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_67_269
timestamp 1698175906
transform 1 0 31472 0 -1 56448
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_67_274
timestamp 1698175906
transform 1 0 32032 0 -1 56448
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_67_281
timestamp 1698175906
transform 1 0 32816 0 -1 56448
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_67_289
timestamp 1698175906
transform 1 0 33712 0 -1 56448
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_67_301
timestamp 1698175906
transform 1 0 35056 0 -1 56448
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_67_305
timestamp 1698175906
transform 1 0 35504 0 -1 56448
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_67_308
timestamp 1698175906
transform 1 0 35840 0 -1 56448
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_67_312
timestamp 1698175906
transform 1 0 36288 0 -1 56448
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_67_321
timestamp 1698175906
transform 1 0 37296 0 -1 56448
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_67_325
timestamp 1698175906
transform 1 0 37744 0 -1 56448
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_67_328
timestamp 1698175906
transform 1 0 38080 0 -1 56448
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_67_332
timestamp 1698175906
transform 1 0 38528 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_67_336
timestamp 1698175906
transform 1 0 38976 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_67_402
timestamp 1698175906
transform 1 0 46368 0 -1 56448
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_67_406
timestamp 1698175906
transform 1 0 46816 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_67_410
timestamp 1698175906
transform 1 0 47264 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_67_412
timestamp 1698175906
transform 1 0 47488 0 -1 56448
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_67_441
timestamp 1698175906
transform 1 0 50736 0 -1 56448
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_67_470
timestamp 1698175906
transform 1 0 53984 0 -1 56448
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_67_504
timestamp 1698175906
transform 1 0 57792 0 -1 56448
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_67_508
timestamp 1698175906
transform 1 0 58240 0 -1 56448
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  input1
timestamp 1698175906
transform 1 0 7504 0 -1 56448
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input2
timestamp 1698175906
transform -1 0 23856 0 -1 56448
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input3
timestamp 1698175906
transform -1 0 26096 0 -1 56448
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input4
timestamp 1698175906
transform -1 0 28896 0 -1 56448
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input5
timestamp 1698175906
transform -1 0 30576 0 -1 56448
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input6
timestamp 1698175906
transform 1 0 32144 0 -1 56448
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input7
timestamp 1698175906
transform 1 0 34384 0 -1 56448
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input8
timestamp 1698175906
transform 1 0 36624 0 -1 56448
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input9
timestamp 1698175906
transform -1 0 40320 0 -1 56448
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  input10
timestamp 1698175906
transform 1 0 16800 0 -1 56448
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  input11
timestamp 1698175906
transform 1 0 18704 0 -1 56448
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input12
timestamp 1698175906
transform 1 0 20944 0 -1 56448
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  input13
timestamp 1698175906
transform 1 0 11984 0 -1 56448
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  input14
timestamp 1698175906
transform 1 0 9744 0 -1 56448
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input15
timestamp 1698175906
transform 1 0 1568 0 1 29792
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input16
timestamp 1698175906
transform 1 0 1568 0 1 48608
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input17
timestamp 1698175906
transform 1 0 1568 0 -1 51744
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input18
timestamp 1698175906
transform 1 0 1568 0 -1 53312
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input19
timestamp 1698175906
transform 1 0 1568 0 -1 54880
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input20
timestamp 1698175906
transform 1 0 1568 0 -1 56448
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input21
timestamp 1698175906
transform -1 0 2912 0 -1 56448
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input22
timestamp 1698175906
transform 1 0 1568 0 1 32928
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  input23
timestamp 1698175906
transform 1 0 1568 0 -1 34496
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input24
timestamp 1698175906
transform 1 0 1568 0 -1 37632
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input25
timestamp 1698175906
transform 1 0 1568 0 1 37632
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input26
timestamp 1698175906
transform 1 0 1568 0 -1 40768
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input27
timestamp 1698175906
transform 1 0 1568 0 1 40768
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input28
timestamp 1698175906
transform 1 0 1568 0 1 42336
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input29
timestamp 1698175906
transform 1 0 1568 0 1 45472
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input30
timestamp 1698175906
transform 1 0 1568 0 -1 47040
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  input31
timestamp 1698175906
transform 1 0 1568 0 1 3136
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  input32
timestamp 1698175906
transform 1 0 1568 0 1 20384
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input33
timestamp 1698175906
transform 1 0 1568 0 1 21952
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input34
timestamp 1698175906
transform 1 0 1568 0 1 23520
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input35
timestamp 1698175906
transform 1 0 1568 0 1 25088
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input36
timestamp 1698175906
transform 1 0 1568 0 -1 28224
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input37
timestamp 1698175906
transform 1 0 2240 0 1 29792
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input38
timestamp 1698175906
transform 1 0 1568 0 -1 4704
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  input39
timestamp 1698175906
transform 1 0 1568 0 -1 6272
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input40
timestamp 1698175906
transform 1 0 1568 0 1 7840
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input41
timestamp 1698175906
transform 1 0 1568 0 1 9408
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input42
timestamp 1698175906
transform 1 0 1568 0 1 10976
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input43
timestamp 1698175906
transform 1 0 1568 0 1 12544
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input44
timestamp 1698175906
transform 1 0 1568 0 -1 15680
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  input45
timestamp 1698175906
transform 1 0 1568 0 -1 17248
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input46
timestamp 1698175906
transform 1 0 1568 0 -1 18816
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input47
timestamp 1698175906
transform -1 0 14896 0 -1 56448
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input48
timestamp 1698175906
transform 1 0 5376 0 -1 56448
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output49 $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 40320 0 -1 56448
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output50
timestamp 1698175906
transform 1 0 43456 0 -1 56448
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output51
timestamp 1698175906
transform 1 0 45584 0 1 54880
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output52
timestamp 1698175906
transform 1 0 47824 0 -1 56448
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output53
timestamp 1698175906
transform 1 0 51072 0 -1 56448
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output54
timestamp 1698175906
transform 1 0 52528 0 1 54880
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output55
timestamp 1698175906
transform 1 0 54880 0 -1 56448
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output56
timestamp 1698175906
transform 1 0 55440 0 1 54880
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_0_Left_68 $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 1344 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_0_Right_0
timestamp 1698175906
transform -1 0 58576 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_1_Left_69
timestamp 1698175906
transform 1 0 1344 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_1_Right_1
timestamp 1698175906
transform -1 0 58576 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_2_Left_70
timestamp 1698175906
transform 1 0 1344 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_2_Right_2
timestamp 1698175906
transform -1 0 58576 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_3_Left_71
timestamp 1698175906
transform 1 0 1344 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_3_Right_3
timestamp 1698175906
transform -1 0 58576 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_4_Left_72
timestamp 1698175906
transform 1 0 1344 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_4_Right_4
timestamp 1698175906
transform -1 0 58576 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_5_Left_73
timestamp 1698175906
transform 1 0 1344 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_5_Right_5
timestamp 1698175906
transform -1 0 58576 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_6_Left_74
timestamp 1698175906
transform 1 0 1344 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_6_Right_6
timestamp 1698175906
transform -1 0 58576 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_7_Left_75
timestamp 1698175906
transform 1 0 1344 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_7_Right_7
timestamp 1698175906
transform -1 0 58576 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_8_Left_76
timestamp 1698175906
transform 1 0 1344 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_8_Right_8
timestamp 1698175906
transform -1 0 58576 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_9_Left_77
timestamp 1698175906
transform 1 0 1344 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_9_Right_9
timestamp 1698175906
transform -1 0 58576 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_10_Left_78
timestamp 1698175906
transform 1 0 1344 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_10_Right_10
timestamp 1698175906
transform -1 0 58576 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_11_Left_79
timestamp 1698175906
transform 1 0 1344 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_11_Right_11
timestamp 1698175906
transform -1 0 58576 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_12_Left_80
timestamp 1698175906
transform 1 0 1344 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_12_Right_12
timestamp 1698175906
transform -1 0 58576 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_13_Left_81
timestamp 1698175906
transform 1 0 1344 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_13_Right_13
timestamp 1698175906
transform -1 0 58576 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_14_Left_82
timestamp 1698175906
transform 1 0 1344 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_14_Right_14
timestamp 1698175906
transform -1 0 58576 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_15_Left_83
timestamp 1698175906
transform 1 0 1344 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_15_Right_15
timestamp 1698175906
transform -1 0 58576 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_16_Left_84
timestamp 1698175906
transform 1 0 1344 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_16_Right_16
timestamp 1698175906
transform -1 0 58576 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_17_Left_85
timestamp 1698175906
transform 1 0 1344 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_17_Right_17
timestamp 1698175906
transform -1 0 58576 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_18_Left_86
timestamp 1698175906
transform 1 0 1344 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_18_Right_18
timestamp 1698175906
transform -1 0 58576 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_19_Left_87
timestamp 1698175906
transform 1 0 1344 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_19_Right_19
timestamp 1698175906
transform -1 0 58576 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_20_Left_88
timestamp 1698175906
transform 1 0 1344 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_20_Right_20
timestamp 1698175906
transform -1 0 58576 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_21_Left_89
timestamp 1698175906
transform 1 0 1344 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_21_Right_21
timestamp 1698175906
transform -1 0 58576 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_22_Left_90
timestamp 1698175906
transform 1 0 1344 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_22_Right_22
timestamp 1698175906
transform -1 0 58576 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_23_Left_91
timestamp 1698175906
transform 1 0 1344 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_23_Right_23
timestamp 1698175906
transform -1 0 58576 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_24_Left_92
timestamp 1698175906
transform 1 0 1344 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_24_Right_24
timestamp 1698175906
transform -1 0 58576 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_25_Left_93
timestamp 1698175906
transform 1 0 1344 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_25_Right_25
timestamp 1698175906
transform -1 0 58576 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_26_Left_94
timestamp 1698175906
transform 1 0 1344 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_26_Right_26
timestamp 1698175906
transform -1 0 58576 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_27_Left_95
timestamp 1698175906
transform 1 0 1344 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_27_Right_27
timestamp 1698175906
transform -1 0 58576 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_28_Left_96
timestamp 1698175906
transform 1 0 1344 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_28_Right_28
timestamp 1698175906
transform -1 0 58576 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_29_Left_97
timestamp 1698175906
transform 1 0 1344 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_29_Right_29
timestamp 1698175906
transform -1 0 58576 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_30_Left_98
timestamp 1698175906
transform 1 0 1344 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_30_Right_30
timestamp 1698175906
transform -1 0 58576 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_31_Left_99
timestamp 1698175906
transform 1 0 1344 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_31_Right_31
timestamp 1698175906
transform -1 0 58576 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_32_Left_100
timestamp 1698175906
transform 1 0 1344 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_32_Right_32
timestamp 1698175906
transform -1 0 58576 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_33_Left_101
timestamp 1698175906
transform 1 0 1344 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_33_Right_33
timestamp 1698175906
transform -1 0 58576 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_34_Left_102
timestamp 1698175906
transform 1 0 1344 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_34_Right_34
timestamp 1698175906
transform -1 0 58576 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_35_Left_103
timestamp 1698175906
transform 1 0 1344 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_35_Right_35
timestamp 1698175906
transform -1 0 58576 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_36_Left_104
timestamp 1698175906
transform 1 0 1344 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_36_Right_36
timestamp 1698175906
transform -1 0 58576 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_37_Left_105
timestamp 1698175906
transform 1 0 1344 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_37_Right_37
timestamp 1698175906
transform -1 0 58576 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_38_Left_106
timestamp 1698175906
transform 1 0 1344 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_38_Right_38
timestamp 1698175906
transform -1 0 58576 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_39_Left_107
timestamp 1698175906
transform 1 0 1344 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_39_Right_39
timestamp 1698175906
transform -1 0 58576 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_40_Left_108
timestamp 1698175906
transform 1 0 1344 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_40_Right_40
timestamp 1698175906
transform -1 0 58576 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_41_Left_109
timestamp 1698175906
transform 1 0 1344 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_41_Right_41
timestamp 1698175906
transform -1 0 58576 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_42_Left_110
timestamp 1698175906
transform 1 0 1344 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_42_Right_42
timestamp 1698175906
transform -1 0 58576 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_43_Left_111
timestamp 1698175906
transform 1 0 1344 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_43_Right_43
timestamp 1698175906
transform -1 0 58576 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_44_Left_112
timestamp 1698175906
transform 1 0 1344 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_44_Right_44
timestamp 1698175906
transform -1 0 58576 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_45_Left_113
timestamp 1698175906
transform 1 0 1344 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_45_Right_45
timestamp 1698175906
transform -1 0 58576 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_46_Left_114
timestamp 1698175906
transform 1 0 1344 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_46_Right_46
timestamp 1698175906
transform -1 0 58576 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_47_Left_115
timestamp 1698175906
transform 1 0 1344 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_47_Right_47
timestamp 1698175906
transform -1 0 58576 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_48_Left_116
timestamp 1698175906
transform 1 0 1344 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_48_Right_48
timestamp 1698175906
transform -1 0 58576 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_49_Left_117
timestamp 1698175906
transform 1 0 1344 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_49_Right_49
timestamp 1698175906
transform -1 0 58576 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_50_Left_118
timestamp 1698175906
transform 1 0 1344 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_50_Right_50
timestamp 1698175906
transform -1 0 58576 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_51_Left_119
timestamp 1698175906
transform 1 0 1344 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_51_Right_51
timestamp 1698175906
transform -1 0 58576 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_52_Left_120
timestamp 1698175906
transform 1 0 1344 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_52_Right_52
timestamp 1698175906
transform -1 0 58576 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_53_Left_121
timestamp 1698175906
transform 1 0 1344 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_53_Right_53
timestamp 1698175906
transform -1 0 58576 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_54_Left_122
timestamp 1698175906
transform 1 0 1344 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_54_Right_54
timestamp 1698175906
transform -1 0 58576 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_55_Left_123
timestamp 1698175906
transform 1 0 1344 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_55_Right_55
timestamp 1698175906
transform -1 0 58576 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_56_Left_124
timestamp 1698175906
transform 1 0 1344 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_56_Right_56
timestamp 1698175906
transform -1 0 58576 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_57_Left_125
timestamp 1698175906
transform 1 0 1344 0 -1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_57_Right_57
timestamp 1698175906
transform -1 0 58576 0 -1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_58_Left_126
timestamp 1698175906
transform 1 0 1344 0 1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_58_Right_58
timestamp 1698175906
transform -1 0 58576 0 1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_59_Left_127
timestamp 1698175906
transform 1 0 1344 0 -1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_59_Right_59
timestamp 1698175906
transform -1 0 58576 0 -1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_60_Left_128
timestamp 1698175906
transform 1 0 1344 0 1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_60_Right_60
timestamp 1698175906
transform -1 0 58576 0 1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_61_Left_129
timestamp 1698175906
transform 1 0 1344 0 -1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_61_Right_61
timestamp 1698175906
transform -1 0 58576 0 -1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_62_Left_130
timestamp 1698175906
transform 1 0 1344 0 1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_62_Right_62
timestamp 1698175906
transform -1 0 58576 0 1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_63_Left_131
timestamp 1698175906
transform 1 0 1344 0 -1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_63_Right_63
timestamp 1698175906
transform -1 0 58576 0 -1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_64_Left_132
timestamp 1698175906
transform 1 0 1344 0 1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_64_Right_64
timestamp 1698175906
transform -1 0 58576 0 1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_65_Left_133
timestamp 1698175906
transform 1 0 1344 0 -1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_65_Right_65
timestamp 1698175906
transform -1 0 58576 0 -1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_66_Left_134
timestamp 1698175906
transform 1 0 1344 0 1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_66_Right_66
timestamp 1698175906
transform -1 0 58576 0 1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_67_Left_135
timestamp 1698175906
transform 1 0 1344 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_67_Right_67
timestamp 1698175906
transform -1 0 58576 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_136 $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 5152 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_137
timestamp 1698175906
transform 1 0 8960 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_138
timestamp 1698175906
transform 1 0 12768 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_139
timestamp 1698175906
transform 1 0 16576 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_140
timestamp 1698175906
transform 1 0 20384 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_141
timestamp 1698175906
transform 1 0 24192 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_142
timestamp 1698175906
transform 1 0 28000 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_143
timestamp 1698175906
transform 1 0 31808 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_144
timestamp 1698175906
transform 1 0 35616 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_145
timestamp 1698175906
transform 1 0 39424 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_146
timestamp 1698175906
transform 1 0 43232 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_147
timestamp 1698175906
transform 1 0 47040 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_148
timestamp 1698175906
transform 1 0 50848 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_149
timestamp 1698175906
transform 1 0 54656 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_1_150
timestamp 1698175906
transform 1 0 9184 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_1_151
timestamp 1698175906
transform 1 0 17024 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_1_152
timestamp 1698175906
transform 1 0 24864 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_1_153
timestamp 1698175906
transform 1 0 32704 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_1_154
timestamp 1698175906
transform 1 0 40544 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_1_155
timestamp 1698175906
transform 1 0 48384 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_1_156
timestamp 1698175906
transform 1 0 56224 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_2_157
timestamp 1698175906
transform 1 0 5264 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_2_158
timestamp 1698175906
transform 1 0 13104 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_2_159
timestamp 1698175906
transform 1 0 20944 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_2_160
timestamp 1698175906
transform 1 0 28784 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_2_161
timestamp 1698175906
transform 1 0 36624 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_2_162
timestamp 1698175906
transform 1 0 44464 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_2_163
timestamp 1698175906
transform 1 0 52304 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_3_164
timestamp 1698175906
transform 1 0 9184 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_3_165
timestamp 1698175906
transform 1 0 17024 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_3_166
timestamp 1698175906
transform 1 0 24864 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_3_167
timestamp 1698175906
transform 1 0 32704 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_3_168
timestamp 1698175906
transform 1 0 40544 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_3_169
timestamp 1698175906
transform 1 0 48384 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_3_170
timestamp 1698175906
transform 1 0 56224 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_4_171
timestamp 1698175906
transform 1 0 5264 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_4_172
timestamp 1698175906
transform 1 0 13104 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_4_173
timestamp 1698175906
transform 1 0 20944 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_4_174
timestamp 1698175906
transform 1 0 28784 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_4_175
timestamp 1698175906
transform 1 0 36624 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_4_176
timestamp 1698175906
transform 1 0 44464 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_4_177
timestamp 1698175906
transform 1 0 52304 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_5_178
timestamp 1698175906
transform 1 0 9184 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_5_179
timestamp 1698175906
transform 1 0 17024 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_5_180
timestamp 1698175906
transform 1 0 24864 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_5_181
timestamp 1698175906
transform 1 0 32704 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_5_182
timestamp 1698175906
transform 1 0 40544 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_5_183
timestamp 1698175906
transform 1 0 48384 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_5_184
timestamp 1698175906
transform 1 0 56224 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_6_185
timestamp 1698175906
transform 1 0 5264 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_6_186
timestamp 1698175906
transform 1 0 13104 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_6_187
timestamp 1698175906
transform 1 0 20944 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_6_188
timestamp 1698175906
transform 1 0 28784 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_6_189
timestamp 1698175906
transform 1 0 36624 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_6_190
timestamp 1698175906
transform 1 0 44464 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_6_191
timestamp 1698175906
transform 1 0 52304 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_7_192
timestamp 1698175906
transform 1 0 9184 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_7_193
timestamp 1698175906
transform 1 0 17024 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_7_194
timestamp 1698175906
transform 1 0 24864 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_7_195
timestamp 1698175906
transform 1 0 32704 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_7_196
timestamp 1698175906
transform 1 0 40544 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_7_197
timestamp 1698175906
transform 1 0 48384 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_7_198
timestamp 1698175906
transform 1 0 56224 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_8_199
timestamp 1698175906
transform 1 0 5264 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_8_200
timestamp 1698175906
transform 1 0 13104 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_8_201
timestamp 1698175906
transform 1 0 20944 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_8_202
timestamp 1698175906
transform 1 0 28784 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_8_203
timestamp 1698175906
transform 1 0 36624 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_8_204
timestamp 1698175906
transform 1 0 44464 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_8_205
timestamp 1698175906
transform 1 0 52304 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_9_206
timestamp 1698175906
transform 1 0 9184 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_9_207
timestamp 1698175906
transform 1 0 17024 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_9_208
timestamp 1698175906
transform 1 0 24864 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_9_209
timestamp 1698175906
transform 1 0 32704 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_9_210
timestamp 1698175906
transform 1 0 40544 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_9_211
timestamp 1698175906
transform 1 0 48384 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_9_212
timestamp 1698175906
transform 1 0 56224 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_10_213
timestamp 1698175906
transform 1 0 5264 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_10_214
timestamp 1698175906
transform 1 0 13104 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_10_215
timestamp 1698175906
transform 1 0 20944 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_10_216
timestamp 1698175906
transform 1 0 28784 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_10_217
timestamp 1698175906
transform 1 0 36624 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_10_218
timestamp 1698175906
transform 1 0 44464 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_10_219
timestamp 1698175906
transform 1 0 52304 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_11_220
timestamp 1698175906
transform 1 0 9184 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_11_221
timestamp 1698175906
transform 1 0 17024 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_11_222
timestamp 1698175906
transform 1 0 24864 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_11_223
timestamp 1698175906
transform 1 0 32704 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_11_224
timestamp 1698175906
transform 1 0 40544 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_11_225
timestamp 1698175906
transform 1 0 48384 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_11_226
timestamp 1698175906
transform 1 0 56224 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_12_227
timestamp 1698175906
transform 1 0 5264 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_12_228
timestamp 1698175906
transform 1 0 13104 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_12_229
timestamp 1698175906
transform 1 0 20944 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_12_230
timestamp 1698175906
transform 1 0 28784 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_12_231
timestamp 1698175906
transform 1 0 36624 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_12_232
timestamp 1698175906
transform 1 0 44464 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_12_233
timestamp 1698175906
transform 1 0 52304 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_13_234
timestamp 1698175906
transform 1 0 9184 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_13_235
timestamp 1698175906
transform 1 0 17024 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_13_236
timestamp 1698175906
transform 1 0 24864 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_13_237
timestamp 1698175906
transform 1 0 32704 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_13_238
timestamp 1698175906
transform 1 0 40544 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_13_239
timestamp 1698175906
transform 1 0 48384 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_13_240
timestamp 1698175906
transform 1 0 56224 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_14_241
timestamp 1698175906
transform 1 0 5264 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_14_242
timestamp 1698175906
transform 1 0 13104 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_14_243
timestamp 1698175906
transform 1 0 20944 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_14_244
timestamp 1698175906
transform 1 0 28784 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_14_245
timestamp 1698175906
transform 1 0 36624 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_14_246
timestamp 1698175906
transform 1 0 44464 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_14_247
timestamp 1698175906
transform 1 0 52304 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_15_248
timestamp 1698175906
transform 1 0 9184 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_15_249
timestamp 1698175906
transform 1 0 17024 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_15_250
timestamp 1698175906
transform 1 0 24864 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_15_251
timestamp 1698175906
transform 1 0 32704 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_15_252
timestamp 1698175906
transform 1 0 40544 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_15_253
timestamp 1698175906
transform 1 0 48384 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_15_254
timestamp 1698175906
transform 1 0 56224 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_16_255
timestamp 1698175906
transform 1 0 5264 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_16_256
timestamp 1698175906
transform 1 0 13104 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_16_257
timestamp 1698175906
transform 1 0 20944 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_16_258
timestamp 1698175906
transform 1 0 28784 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_16_259
timestamp 1698175906
transform 1 0 36624 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_16_260
timestamp 1698175906
transform 1 0 44464 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_16_261
timestamp 1698175906
transform 1 0 52304 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_17_262
timestamp 1698175906
transform 1 0 9184 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_17_263
timestamp 1698175906
transform 1 0 17024 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_17_264
timestamp 1698175906
transform 1 0 24864 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_17_265
timestamp 1698175906
transform 1 0 32704 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_17_266
timestamp 1698175906
transform 1 0 40544 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_17_267
timestamp 1698175906
transform 1 0 48384 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_17_268
timestamp 1698175906
transform 1 0 56224 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_18_269
timestamp 1698175906
transform 1 0 5264 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_18_270
timestamp 1698175906
transform 1 0 13104 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_18_271
timestamp 1698175906
transform 1 0 20944 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_18_272
timestamp 1698175906
transform 1 0 28784 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_18_273
timestamp 1698175906
transform 1 0 36624 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_18_274
timestamp 1698175906
transform 1 0 44464 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_18_275
timestamp 1698175906
transform 1 0 52304 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_19_276
timestamp 1698175906
transform 1 0 9184 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_19_277
timestamp 1698175906
transform 1 0 17024 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_19_278
timestamp 1698175906
transform 1 0 24864 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_19_279
timestamp 1698175906
transform 1 0 32704 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_19_280
timestamp 1698175906
transform 1 0 40544 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_19_281
timestamp 1698175906
transform 1 0 48384 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_19_282
timestamp 1698175906
transform 1 0 56224 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_20_283
timestamp 1698175906
transform 1 0 5264 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_20_284
timestamp 1698175906
transform 1 0 13104 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_20_285
timestamp 1698175906
transform 1 0 20944 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_20_286
timestamp 1698175906
transform 1 0 28784 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_20_287
timestamp 1698175906
transform 1 0 36624 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_20_288
timestamp 1698175906
transform 1 0 44464 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_20_289
timestamp 1698175906
transform 1 0 52304 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_21_290
timestamp 1698175906
transform 1 0 9184 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_21_291
timestamp 1698175906
transform 1 0 17024 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_21_292
timestamp 1698175906
transform 1 0 24864 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_21_293
timestamp 1698175906
transform 1 0 32704 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_21_294
timestamp 1698175906
transform 1 0 40544 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_21_295
timestamp 1698175906
transform 1 0 48384 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_21_296
timestamp 1698175906
transform 1 0 56224 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_22_297
timestamp 1698175906
transform 1 0 5264 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_22_298
timestamp 1698175906
transform 1 0 13104 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_22_299
timestamp 1698175906
transform 1 0 20944 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_22_300
timestamp 1698175906
transform 1 0 28784 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_22_301
timestamp 1698175906
transform 1 0 36624 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_22_302
timestamp 1698175906
transform 1 0 44464 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_22_303
timestamp 1698175906
transform 1 0 52304 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_23_304
timestamp 1698175906
transform 1 0 9184 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_23_305
timestamp 1698175906
transform 1 0 17024 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_23_306
timestamp 1698175906
transform 1 0 24864 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_23_307
timestamp 1698175906
transform 1 0 32704 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_23_308
timestamp 1698175906
transform 1 0 40544 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_23_309
timestamp 1698175906
transform 1 0 48384 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_23_310
timestamp 1698175906
transform 1 0 56224 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_24_311
timestamp 1698175906
transform 1 0 5264 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_24_312
timestamp 1698175906
transform 1 0 13104 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_24_313
timestamp 1698175906
transform 1 0 20944 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_24_314
timestamp 1698175906
transform 1 0 28784 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_24_315
timestamp 1698175906
transform 1 0 36624 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_24_316
timestamp 1698175906
transform 1 0 44464 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_24_317
timestamp 1698175906
transform 1 0 52304 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_25_318
timestamp 1698175906
transform 1 0 9184 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_25_319
timestamp 1698175906
transform 1 0 17024 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_25_320
timestamp 1698175906
transform 1 0 24864 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_25_321
timestamp 1698175906
transform 1 0 32704 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_25_322
timestamp 1698175906
transform 1 0 40544 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_25_323
timestamp 1698175906
transform 1 0 48384 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_25_324
timestamp 1698175906
transform 1 0 56224 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_26_325
timestamp 1698175906
transform 1 0 5264 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_26_326
timestamp 1698175906
transform 1 0 13104 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_26_327
timestamp 1698175906
transform 1 0 20944 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_26_328
timestamp 1698175906
transform 1 0 28784 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_26_329
timestamp 1698175906
transform 1 0 36624 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_26_330
timestamp 1698175906
transform 1 0 44464 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_26_331
timestamp 1698175906
transform 1 0 52304 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_27_332
timestamp 1698175906
transform 1 0 9184 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_27_333
timestamp 1698175906
transform 1 0 17024 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_27_334
timestamp 1698175906
transform 1 0 24864 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_27_335
timestamp 1698175906
transform 1 0 32704 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_27_336
timestamp 1698175906
transform 1 0 40544 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_27_337
timestamp 1698175906
transform 1 0 48384 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_27_338
timestamp 1698175906
transform 1 0 56224 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_28_339
timestamp 1698175906
transform 1 0 5264 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_28_340
timestamp 1698175906
transform 1 0 13104 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_28_341
timestamp 1698175906
transform 1 0 20944 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_28_342
timestamp 1698175906
transform 1 0 28784 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_28_343
timestamp 1698175906
transform 1 0 36624 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_28_344
timestamp 1698175906
transform 1 0 44464 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_28_345
timestamp 1698175906
transform 1 0 52304 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_29_346
timestamp 1698175906
transform 1 0 9184 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_29_347
timestamp 1698175906
transform 1 0 17024 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_29_348
timestamp 1698175906
transform 1 0 24864 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_29_349
timestamp 1698175906
transform 1 0 32704 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_29_350
timestamp 1698175906
transform 1 0 40544 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_29_351
timestamp 1698175906
transform 1 0 48384 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_29_352
timestamp 1698175906
transform 1 0 56224 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_30_353
timestamp 1698175906
transform 1 0 5264 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_30_354
timestamp 1698175906
transform 1 0 13104 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_30_355
timestamp 1698175906
transform 1 0 20944 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_30_356
timestamp 1698175906
transform 1 0 28784 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_30_357
timestamp 1698175906
transform 1 0 36624 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_30_358
timestamp 1698175906
transform 1 0 44464 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_30_359
timestamp 1698175906
transform 1 0 52304 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_31_360
timestamp 1698175906
transform 1 0 9184 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_31_361
timestamp 1698175906
transform 1 0 17024 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_31_362
timestamp 1698175906
transform 1 0 24864 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_31_363
timestamp 1698175906
transform 1 0 32704 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_31_364
timestamp 1698175906
transform 1 0 40544 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_31_365
timestamp 1698175906
transform 1 0 48384 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_31_366
timestamp 1698175906
transform 1 0 56224 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_32_367
timestamp 1698175906
transform 1 0 5264 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_32_368
timestamp 1698175906
transform 1 0 13104 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_32_369
timestamp 1698175906
transform 1 0 20944 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_32_370
timestamp 1698175906
transform 1 0 28784 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_32_371
timestamp 1698175906
transform 1 0 36624 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_32_372
timestamp 1698175906
transform 1 0 44464 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_32_373
timestamp 1698175906
transform 1 0 52304 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_33_374
timestamp 1698175906
transform 1 0 9184 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_33_375
timestamp 1698175906
transform 1 0 17024 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_33_376
timestamp 1698175906
transform 1 0 24864 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_33_377
timestamp 1698175906
transform 1 0 32704 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_33_378
timestamp 1698175906
transform 1 0 40544 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_33_379
timestamp 1698175906
transform 1 0 48384 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_33_380
timestamp 1698175906
transform 1 0 56224 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_34_381
timestamp 1698175906
transform 1 0 5264 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_34_382
timestamp 1698175906
transform 1 0 13104 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_34_383
timestamp 1698175906
transform 1 0 20944 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_34_384
timestamp 1698175906
transform 1 0 28784 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_34_385
timestamp 1698175906
transform 1 0 36624 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_34_386
timestamp 1698175906
transform 1 0 44464 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_34_387
timestamp 1698175906
transform 1 0 52304 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_35_388
timestamp 1698175906
transform 1 0 9184 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_35_389
timestamp 1698175906
transform 1 0 17024 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_35_390
timestamp 1698175906
transform 1 0 24864 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_35_391
timestamp 1698175906
transform 1 0 32704 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_35_392
timestamp 1698175906
transform 1 0 40544 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_35_393
timestamp 1698175906
transform 1 0 48384 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_35_394
timestamp 1698175906
transform 1 0 56224 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_36_395
timestamp 1698175906
transform 1 0 5264 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_36_396
timestamp 1698175906
transform 1 0 13104 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_36_397
timestamp 1698175906
transform 1 0 20944 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_36_398
timestamp 1698175906
transform 1 0 28784 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_36_399
timestamp 1698175906
transform 1 0 36624 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_36_400
timestamp 1698175906
transform 1 0 44464 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_36_401
timestamp 1698175906
transform 1 0 52304 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_37_402
timestamp 1698175906
transform 1 0 9184 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_37_403
timestamp 1698175906
transform 1 0 17024 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_37_404
timestamp 1698175906
transform 1 0 24864 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_37_405
timestamp 1698175906
transform 1 0 32704 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_37_406
timestamp 1698175906
transform 1 0 40544 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_37_407
timestamp 1698175906
transform 1 0 48384 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_37_408
timestamp 1698175906
transform 1 0 56224 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_38_409
timestamp 1698175906
transform 1 0 5264 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_38_410
timestamp 1698175906
transform 1 0 13104 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_38_411
timestamp 1698175906
transform 1 0 20944 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_38_412
timestamp 1698175906
transform 1 0 28784 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_38_413
timestamp 1698175906
transform 1 0 36624 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_38_414
timestamp 1698175906
transform 1 0 44464 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_38_415
timestamp 1698175906
transform 1 0 52304 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_39_416
timestamp 1698175906
transform 1 0 9184 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_39_417
timestamp 1698175906
transform 1 0 17024 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_39_418
timestamp 1698175906
transform 1 0 24864 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_39_419
timestamp 1698175906
transform 1 0 32704 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_39_420
timestamp 1698175906
transform 1 0 40544 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_39_421
timestamp 1698175906
transform 1 0 48384 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_39_422
timestamp 1698175906
transform 1 0 56224 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_40_423
timestamp 1698175906
transform 1 0 5264 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_40_424
timestamp 1698175906
transform 1 0 13104 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_40_425
timestamp 1698175906
transform 1 0 20944 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_40_426
timestamp 1698175906
transform 1 0 28784 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_40_427
timestamp 1698175906
transform 1 0 36624 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_40_428
timestamp 1698175906
transform 1 0 44464 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_40_429
timestamp 1698175906
transform 1 0 52304 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_41_430
timestamp 1698175906
transform 1 0 9184 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_41_431
timestamp 1698175906
transform 1 0 17024 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_41_432
timestamp 1698175906
transform 1 0 24864 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_41_433
timestamp 1698175906
transform 1 0 32704 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_41_434
timestamp 1698175906
transform 1 0 40544 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_41_435
timestamp 1698175906
transform 1 0 48384 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_41_436
timestamp 1698175906
transform 1 0 56224 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_42_437
timestamp 1698175906
transform 1 0 5264 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_42_438
timestamp 1698175906
transform 1 0 13104 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_42_439
timestamp 1698175906
transform 1 0 20944 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_42_440
timestamp 1698175906
transform 1 0 28784 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_42_441
timestamp 1698175906
transform 1 0 36624 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_42_442
timestamp 1698175906
transform 1 0 44464 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_42_443
timestamp 1698175906
transform 1 0 52304 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_43_444
timestamp 1698175906
transform 1 0 9184 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_43_445
timestamp 1698175906
transform 1 0 17024 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_43_446
timestamp 1698175906
transform 1 0 24864 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_43_447
timestamp 1698175906
transform 1 0 32704 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_43_448
timestamp 1698175906
transform 1 0 40544 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_43_449
timestamp 1698175906
transform 1 0 48384 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_43_450
timestamp 1698175906
transform 1 0 56224 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_44_451
timestamp 1698175906
transform 1 0 5264 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_44_452
timestamp 1698175906
transform 1 0 13104 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_44_453
timestamp 1698175906
transform 1 0 20944 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_44_454
timestamp 1698175906
transform 1 0 28784 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_44_455
timestamp 1698175906
transform 1 0 36624 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_44_456
timestamp 1698175906
transform 1 0 44464 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_44_457
timestamp 1698175906
transform 1 0 52304 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_45_458
timestamp 1698175906
transform 1 0 9184 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_45_459
timestamp 1698175906
transform 1 0 17024 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_45_460
timestamp 1698175906
transform 1 0 24864 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_45_461
timestamp 1698175906
transform 1 0 32704 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_45_462
timestamp 1698175906
transform 1 0 40544 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_45_463
timestamp 1698175906
transform 1 0 48384 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_45_464
timestamp 1698175906
transform 1 0 56224 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_46_465
timestamp 1698175906
transform 1 0 5264 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_46_466
timestamp 1698175906
transform 1 0 13104 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_46_467
timestamp 1698175906
transform 1 0 20944 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_46_468
timestamp 1698175906
transform 1 0 28784 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_46_469
timestamp 1698175906
transform 1 0 36624 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_46_470
timestamp 1698175906
transform 1 0 44464 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_46_471
timestamp 1698175906
transform 1 0 52304 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_47_472
timestamp 1698175906
transform 1 0 9184 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_47_473
timestamp 1698175906
transform 1 0 17024 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_47_474
timestamp 1698175906
transform 1 0 24864 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_47_475
timestamp 1698175906
transform 1 0 32704 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_47_476
timestamp 1698175906
transform 1 0 40544 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_47_477
timestamp 1698175906
transform 1 0 48384 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_47_478
timestamp 1698175906
transform 1 0 56224 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_48_479
timestamp 1698175906
transform 1 0 5264 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_48_480
timestamp 1698175906
transform 1 0 13104 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_48_481
timestamp 1698175906
transform 1 0 20944 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_48_482
timestamp 1698175906
transform 1 0 28784 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_48_483
timestamp 1698175906
transform 1 0 36624 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_48_484
timestamp 1698175906
transform 1 0 44464 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_48_485
timestamp 1698175906
transform 1 0 52304 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_49_486
timestamp 1698175906
transform 1 0 9184 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_49_487
timestamp 1698175906
transform 1 0 17024 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_49_488
timestamp 1698175906
transform 1 0 24864 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_49_489
timestamp 1698175906
transform 1 0 32704 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_49_490
timestamp 1698175906
transform 1 0 40544 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_49_491
timestamp 1698175906
transform 1 0 48384 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_49_492
timestamp 1698175906
transform 1 0 56224 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_50_493
timestamp 1698175906
transform 1 0 5264 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_50_494
timestamp 1698175906
transform 1 0 13104 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_50_495
timestamp 1698175906
transform 1 0 20944 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_50_496
timestamp 1698175906
transform 1 0 28784 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_50_497
timestamp 1698175906
transform 1 0 36624 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_50_498
timestamp 1698175906
transform 1 0 44464 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_50_499
timestamp 1698175906
transform 1 0 52304 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_51_500
timestamp 1698175906
transform 1 0 9184 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_51_501
timestamp 1698175906
transform 1 0 17024 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_51_502
timestamp 1698175906
transform 1 0 24864 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_51_503
timestamp 1698175906
transform 1 0 32704 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_51_504
timestamp 1698175906
transform 1 0 40544 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_51_505
timestamp 1698175906
transform 1 0 48384 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_51_506
timestamp 1698175906
transform 1 0 56224 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_52_507
timestamp 1698175906
transform 1 0 5264 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_52_508
timestamp 1698175906
transform 1 0 13104 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_52_509
timestamp 1698175906
transform 1 0 20944 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_52_510
timestamp 1698175906
transform 1 0 28784 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_52_511
timestamp 1698175906
transform 1 0 36624 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_52_512
timestamp 1698175906
transform 1 0 44464 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_52_513
timestamp 1698175906
transform 1 0 52304 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_53_514
timestamp 1698175906
transform 1 0 9184 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_53_515
timestamp 1698175906
transform 1 0 17024 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_53_516
timestamp 1698175906
transform 1 0 24864 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_53_517
timestamp 1698175906
transform 1 0 32704 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_53_518
timestamp 1698175906
transform 1 0 40544 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_53_519
timestamp 1698175906
transform 1 0 48384 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_53_520
timestamp 1698175906
transform 1 0 56224 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_54_521
timestamp 1698175906
transform 1 0 5264 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_54_522
timestamp 1698175906
transform 1 0 13104 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_54_523
timestamp 1698175906
transform 1 0 20944 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_54_524
timestamp 1698175906
transform 1 0 28784 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_54_525
timestamp 1698175906
transform 1 0 36624 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_54_526
timestamp 1698175906
transform 1 0 44464 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_54_527
timestamp 1698175906
transform 1 0 52304 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_55_528
timestamp 1698175906
transform 1 0 9184 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_55_529
timestamp 1698175906
transform 1 0 17024 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_55_530
timestamp 1698175906
transform 1 0 24864 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_55_531
timestamp 1698175906
transform 1 0 32704 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_55_532
timestamp 1698175906
transform 1 0 40544 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_55_533
timestamp 1698175906
transform 1 0 48384 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_55_534
timestamp 1698175906
transform 1 0 56224 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_56_535
timestamp 1698175906
transform 1 0 5264 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_56_536
timestamp 1698175906
transform 1 0 13104 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_56_537
timestamp 1698175906
transform 1 0 20944 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_56_538
timestamp 1698175906
transform 1 0 28784 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_56_539
timestamp 1698175906
transform 1 0 36624 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_56_540
timestamp 1698175906
transform 1 0 44464 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_56_541
timestamp 1698175906
transform 1 0 52304 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_57_542
timestamp 1698175906
transform 1 0 9184 0 -1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_57_543
timestamp 1698175906
transform 1 0 17024 0 -1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_57_544
timestamp 1698175906
transform 1 0 24864 0 -1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_57_545
timestamp 1698175906
transform 1 0 32704 0 -1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_57_546
timestamp 1698175906
transform 1 0 40544 0 -1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_57_547
timestamp 1698175906
transform 1 0 48384 0 -1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_57_548
timestamp 1698175906
transform 1 0 56224 0 -1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_58_549
timestamp 1698175906
transform 1 0 5264 0 1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_58_550
timestamp 1698175906
transform 1 0 13104 0 1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_58_551
timestamp 1698175906
transform 1 0 20944 0 1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_58_552
timestamp 1698175906
transform 1 0 28784 0 1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_58_553
timestamp 1698175906
transform 1 0 36624 0 1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_58_554
timestamp 1698175906
transform 1 0 44464 0 1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_58_555
timestamp 1698175906
transform 1 0 52304 0 1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_59_556
timestamp 1698175906
transform 1 0 9184 0 -1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_59_557
timestamp 1698175906
transform 1 0 17024 0 -1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_59_558
timestamp 1698175906
transform 1 0 24864 0 -1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_59_559
timestamp 1698175906
transform 1 0 32704 0 -1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_59_560
timestamp 1698175906
transform 1 0 40544 0 -1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_59_561
timestamp 1698175906
transform 1 0 48384 0 -1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_59_562
timestamp 1698175906
transform 1 0 56224 0 -1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_60_563
timestamp 1698175906
transform 1 0 5264 0 1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_60_564
timestamp 1698175906
transform 1 0 13104 0 1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_60_565
timestamp 1698175906
transform 1 0 20944 0 1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_60_566
timestamp 1698175906
transform 1 0 28784 0 1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_60_567
timestamp 1698175906
transform 1 0 36624 0 1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_60_568
timestamp 1698175906
transform 1 0 44464 0 1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_60_569
timestamp 1698175906
transform 1 0 52304 0 1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_61_570
timestamp 1698175906
transform 1 0 9184 0 -1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_61_571
timestamp 1698175906
transform 1 0 17024 0 -1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_61_572
timestamp 1698175906
transform 1 0 24864 0 -1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_61_573
timestamp 1698175906
transform 1 0 32704 0 -1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_61_574
timestamp 1698175906
transform 1 0 40544 0 -1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_61_575
timestamp 1698175906
transform 1 0 48384 0 -1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_61_576
timestamp 1698175906
transform 1 0 56224 0 -1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_62_577
timestamp 1698175906
transform 1 0 5264 0 1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_62_578
timestamp 1698175906
transform 1 0 13104 0 1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_62_579
timestamp 1698175906
transform 1 0 20944 0 1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_62_580
timestamp 1698175906
transform 1 0 28784 0 1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_62_581
timestamp 1698175906
transform 1 0 36624 0 1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_62_582
timestamp 1698175906
transform 1 0 44464 0 1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_62_583
timestamp 1698175906
transform 1 0 52304 0 1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_63_584
timestamp 1698175906
transform 1 0 9184 0 -1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_63_585
timestamp 1698175906
transform 1 0 17024 0 -1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_63_586
timestamp 1698175906
transform 1 0 24864 0 -1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_63_587
timestamp 1698175906
transform 1 0 32704 0 -1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_63_588
timestamp 1698175906
transform 1 0 40544 0 -1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_63_589
timestamp 1698175906
transform 1 0 48384 0 -1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_63_590
timestamp 1698175906
transform 1 0 56224 0 -1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_64_591
timestamp 1698175906
transform 1 0 5264 0 1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_64_592
timestamp 1698175906
transform 1 0 13104 0 1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_64_593
timestamp 1698175906
transform 1 0 20944 0 1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_64_594
timestamp 1698175906
transform 1 0 28784 0 1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_64_595
timestamp 1698175906
transform 1 0 36624 0 1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_64_596
timestamp 1698175906
transform 1 0 44464 0 1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_64_597
timestamp 1698175906
transform 1 0 52304 0 1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_65_598
timestamp 1698175906
transform 1 0 9184 0 -1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_65_599
timestamp 1698175906
transform 1 0 17024 0 -1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_65_600
timestamp 1698175906
transform 1 0 24864 0 -1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_65_601
timestamp 1698175906
transform 1 0 32704 0 -1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_65_602
timestamp 1698175906
transform 1 0 40544 0 -1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_65_603
timestamp 1698175906
transform 1 0 48384 0 -1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_65_604
timestamp 1698175906
transform 1 0 56224 0 -1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_66_605
timestamp 1698175906
transform 1 0 5264 0 1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_66_606
timestamp 1698175906
transform 1 0 13104 0 1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_66_607
timestamp 1698175906
transform 1 0 20944 0 1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_66_608
timestamp 1698175906
transform 1 0 28784 0 1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_66_609
timestamp 1698175906
transform 1 0 36624 0 1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_66_610
timestamp 1698175906
transform 1 0 44464 0 1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_66_611
timestamp 1698175906
transform 1 0 52304 0 1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_67_612
timestamp 1698175906
transform 1 0 5152 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_67_613
timestamp 1698175906
transform 1 0 8960 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_67_614
timestamp 1698175906
transform 1 0 12768 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_67_615
timestamp 1698175906
transform 1 0 16576 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_67_616
timestamp 1698175906
transform 1 0 20384 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_67_617
timestamp 1698175906
transform 1 0 24192 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_67_618
timestamp 1698175906
transform 1 0 28000 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_67_619
timestamp 1698175906
transform 1 0 31808 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_67_620
timestamp 1698175906
transform 1 0 35616 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_67_621
timestamp 1698175906
transform 1 0 39424 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_67_622
timestamp 1698175906
transform 1 0 43232 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_67_623
timestamp 1698175906
transform 1 0 47040 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_67_624
timestamp 1698175906
transform 1 0 50848 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_67_625
timestamp 1698175906
transform 1 0 54656 0 -1 56448
box -86 -86 310 870
<< labels >>
flabel metal2 s 7392 59200 7504 60000 0 FreeSans 448 90 0 0 WEb_raw
port 0 nsew signal input
flabel metal2 s 23072 59200 23184 60000 0 FreeSans 448 90 0 0 bus_in[0]
port 1 nsew signal input
flabel metal2 s 25312 59200 25424 60000 0 FreeSans 448 90 0 0 bus_in[1]
port 2 nsew signal input
flabel metal2 s 27552 59200 27664 60000 0 FreeSans 448 90 0 0 bus_in[2]
port 3 nsew signal input
flabel metal2 s 29792 59200 29904 60000 0 FreeSans 448 90 0 0 bus_in[3]
port 4 nsew signal input
flabel metal2 s 32032 59200 32144 60000 0 FreeSans 448 90 0 0 bus_in[4]
port 5 nsew signal input
flabel metal2 s 34272 59200 34384 60000 0 FreeSans 448 90 0 0 bus_in[5]
port 6 nsew signal input
flabel metal2 s 36512 59200 36624 60000 0 FreeSans 448 90 0 0 bus_in[6]
port 7 nsew signal input
flabel metal2 s 38752 59200 38864 60000 0 FreeSans 448 90 0 0 bus_in[7]
port 8 nsew signal input
flabel metal2 s 40992 59200 41104 60000 0 FreeSans 448 90 0 0 bus_out[0]
port 9 nsew signal tristate
flabel metal2 s 43232 59200 43344 60000 0 FreeSans 448 90 0 0 bus_out[1]
port 10 nsew signal tristate
flabel metal2 s 45472 59200 45584 60000 0 FreeSans 448 90 0 0 bus_out[2]
port 11 nsew signal tristate
flabel metal2 s 47712 59200 47824 60000 0 FreeSans 448 90 0 0 bus_out[3]
port 12 nsew signal tristate
flabel metal2 s 49952 59200 50064 60000 0 FreeSans 448 90 0 0 bus_out[4]
port 13 nsew signal tristate
flabel metal2 s 52192 59200 52304 60000 0 FreeSans 448 90 0 0 bus_out[5]
port 14 nsew signal tristate
flabel metal2 s 54432 59200 54544 60000 0 FreeSans 448 90 0 0 bus_out[6]
port 15 nsew signal tristate
flabel metal2 s 56672 59200 56784 60000 0 FreeSans 448 90 0 0 bus_out[7]
port 16 nsew signal tristate
flabel metal2 s 16352 59200 16464 60000 0 FreeSans 448 90 0 0 cs_port[0]
port 17 nsew signal input
flabel metal2 s 18592 59200 18704 60000 0 FreeSans 448 90 0 0 cs_port[1]
port 18 nsew signal input
flabel metal2 s 20832 59200 20944 60000 0 FreeSans 448 90 0 0 cs_port[2]
port 19 nsew signal input
flabel metal2 s 11872 59200 11984 60000 0 FreeSans 448 90 0 0 le_hi_act
port 20 nsew signal input
flabel metal2 s 9632 59200 9744 60000 0 FreeSans 448 90 0 0 le_lo_act
port 21 nsew signal input
flabel metal3 s 0 30688 800 30800 0 FreeSans 448 0 0 0 ram_end[0]
port 22 nsew signal input
flabel metal3 s 0 48608 800 48720 0 FreeSans 448 0 0 0 ram_end[10]
port 23 nsew signal input
flabel metal3 s 0 50400 800 50512 0 FreeSans 448 0 0 0 ram_end[11]
port 24 nsew signal input
flabel metal3 s 0 52192 800 52304 0 FreeSans 448 0 0 0 ram_end[12]
port 25 nsew signal input
flabel metal3 s 0 53984 800 54096 0 FreeSans 448 0 0 0 ram_end[13]
port 26 nsew signal input
flabel metal3 s 0 55776 800 55888 0 FreeSans 448 0 0 0 ram_end[14]
port 27 nsew signal input
flabel metal3 s 0 57568 800 57680 0 FreeSans 448 0 0 0 ram_end[15]
port 28 nsew signal input
flabel metal3 s 0 32480 800 32592 0 FreeSans 448 0 0 0 ram_end[1]
port 29 nsew signal input
flabel metal3 s 0 34272 800 34384 0 FreeSans 448 0 0 0 ram_end[2]
port 30 nsew signal input
flabel metal3 s 0 36064 800 36176 0 FreeSans 448 0 0 0 ram_end[3]
port 31 nsew signal input
flabel metal3 s 0 37856 800 37968 0 FreeSans 448 0 0 0 ram_end[4]
port 32 nsew signal input
flabel metal3 s 0 39648 800 39760 0 FreeSans 448 0 0 0 ram_end[5]
port 33 nsew signal input
flabel metal3 s 0 41440 800 41552 0 FreeSans 448 0 0 0 ram_end[6]
port 34 nsew signal input
flabel metal3 s 0 43232 800 43344 0 FreeSans 448 0 0 0 ram_end[7]
port 35 nsew signal input
flabel metal3 s 0 45024 800 45136 0 FreeSans 448 0 0 0 ram_end[8]
port 36 nsew signal input
flabel metal3 s 0 46816 800 46928 0 FreeSans 448 0 0 0 ram_end[9]
port 37 nsew signal input
flabel metal3 s 0 2016 800 2128 0 FreeSans 448 0 0 0 ram_start[0]
port 38 nsew signal input
flabel metal3 s 0 19936 800 20048 0 FreeSans 448 0 0 0 ram_start[10]
port 39 nsew signal input
flabel metal3 s 0 21728 800 21840 0 FreeSans 448 0 0 0 ram_start[11]
port 40 nsew signal input
flabel metal3 s 0 23520 800 23632 0 FreeSans 448 0 0 0 ram_start[12]
port 41 nsew signal input
flabel metal3 s 0 25312 800 25424 0 FreeSans 448 0 0 0 ram_start[13]
port 42 nsew signal input
flabel metal3 s 0 27104 800 27216 0 FreeSans 448 0 0 0 ram_start[14]
port 43 nsew signal input
flabel metal3 s 0 28896 800 29008 0 FreeSans 448 0 0 0 ram_start[15]
port 44 nsew signal input
flabel metal3 s 0 3808 800 3920 0 FreeSans 448 0 0 0 ram_start[1]
port 45 nsew signal input
flabel metal3 s 0 5600 800 5712 0 FreeSans 448 0 0 0 ram_start[2]
port 46 nsew signal input
flabel metal3 s 0 7392 800 7504 0 FreeSans 448 0 0 0 ram_start[3]
port 47 nsew signal input
flabel metal3 s 0 9184 800 9296 0 FreeSans 448 0 0 0 ram_start[4]
port 48 nsew signal input
flabel metal3 s 0 10976 800 11088 0 FreeSans 448 0 0 0 ram_start[5]
port 49 nsew signal input
flabel metal3 s 0 12768 800 12880 0 FreeSans 448 0 0 0 ram_start[6]
port 50 nsew signal input
flabel metal3 s 0 14560 800 14672 0 FreeSans 448 0 0 0 ram_start[7]
port 51 nsew signal input
flabel metal3 s 0 16352 800 16464 0 FreeSans 448 0 0 0 ram_start[8]
port 52 nsew signal input
flabel metal3 s 0 18144 800 18256 0 FreeSans 448 0 0 0 ram_start[9]
port 53 nsew signal input
flabel metal2 s 14112 59200 14224 60000 0 FreeSans 448 90 0 0 rom_enabled
port 54 nsew signal input
flabel metal2 s 5152 59200 5264 60000 0 FreeSans 448 90 0 0 rst
port 55 nsew signal input
flabel metal4 s 4448 3076 4768 56508 0 FreeSans 1280 90 0 0 vdd
port 56 nsew power bidirectional
flabel metal4 s 35168 3076 35488 56508 0 FreeSans 1280 90 0 0 vdd
port 56 nsew power bidirectional
flabel metal4 s 19808 3076 20128 56508 0 FreeSans 1280 90 0 0 vss
port 57 nsew ground bidirectional
flabel metal4 s 50528 3076 50848 56508 0 FreeSans 1280 90 0 0 vss
port 57 nsew ground bidirectional
flabel metal2 s 2912 59200 3024 60000 0 FreeSans 448 90 0 0 wb_clk_i
port 58 nsew signal input
rlabel metal1 29960 55664 29960 55664 0 vdd
rlabel metal1 29960 56448 29960 56448 0 vss
rlabel metal2 7448 57778 7448 57778 0 WEb_raw
rlabel metal3 7336 49896 7336 49896 0 _0000_
rlabel metal2 3864 51296 3864 51296 0 _0001_
rlabel metal3 9352 52920 9352 52920 0 _0002_
rlabel metal2 11928 51576 11928 51576 0 _0003_
rlabel metal2 37800 41216 37800 41216 0 _0004_
rlabel metal3 35560 40264 35560 40264 0 _0005_
rlabel metal3 37016 38920 37016 38920 0 _0006_
rlabel metal2 34664 43848 34664 43848 0 _0007_
rlabel metal2 21784 52136 21784 52136 0 _0008_
rlabel metal2 24920 53928 24920 53928 0 _0009_
rlabel metal3 22120 53704 22120 53704 0 _0010_
rlabel metal2 26488 50960 26488 50960 0 _0011_
rlabel metal2 41272 47096 41272 47096 0 _0012_
rlabel metal2 40488 42560 40488 42560 0 _0013_
rlabel metal2 39368 43848 39368 43848 0 _0014_
rlabel metal2 42392 45248 42392 45248 0 _0015_
rlabel metal2 29960 54936 29960 54936 0 _0016_
rlabel metal2 30184 52528 30184 52528 0 _0017_
rlabel metal2 34328 54936 34328 54936 0 _0018_
rlabel metal2 34216 52696 34216 52696 0 _0019_
rlabel metal2 37912 50960 37912 50960 0 _0020_
rlabel metal2 41384 52472 41384 52472 0 _0021_
rlabel metal2 42056 50848 42056 50848 0 _0022_
rlabel metal2 41048 54936 41048 54936 0 _0023_
rlabel metal2 14840 54936 14840 54936 0 _0024_
rlabel metal2 13944 51576 13944 51576 0 _0025_
rlabel metal2 17640 54768 17640 54768 0 _0026_
rlabel metal2 19992 52528 19992 52528 0 _0027_
rlabel metal2 33320 46872 33320 46872 0 _0028_
rlabel metal2 35672 49392 35672 49392 0 _0029_
rlabel metal3 35952 46760 35952 46760 0 _0030_
rlabel metal2 31416 49056 31416 49056 0 _0031_
rlabel metal2 25368 49056 25368 49056 0 _0032_
rlabel metal2 37464 52416 37464 52416 0 _0033_
rlabel metal3 40768 52024 40768 52024 0 _0034_
rlabel metal2 38696 51912 38696 51912 0 _0035_
rlabel metal2 37464 30184 37464 30184 0 _0036_
rlabel metal2 33152 36456 33152 36456 0 _0037_
rlabel metal2 35224 32928 35224 32928 0 _0038_
rlabel metal2 39144 35224 39144 35224 0 _0039_
rlabel metal2 34328 39872 34328 39872 0 _0040_
rlabel metal2 38920 33824 38920 33824 0 _0041_
rlabel metal2 15736 46480 15736 46480 0 _0042_
rlabel metal2 6664 47096 6664 47096 0 _0043_
rlabel metal3 5600 40488 5600 40488 0 _0044_
rlabel metal2 7336 48160 7336 48160 0 _0045_
rlabel metal2 9800 43008 9800 43008 0 _0046_
rlabel metal2 8344 47936 8344 47936 0 _0047_
rlabel metal2 12152 45808 12152 45808 0 _0048_
rlabel metal2 2520 47488 2520 47488 0 _0049_
rlabel metal3 6384 46760 6384 46760 0 _0050_
rlabel metal2 10248 45024 10248 45024 0 _0051_
rlabel metal2 13944 47824 13944 47824 0 _0052_
rlabel metal3 20664 40600 20664 40600 0 _0053_
rlabel metal2 26040 45920 26040 45920 0 _0054_
rlabel metal2 39592 34440 39592 34440 0 _0055_
rlabel metal2 39256 35840 39256 35840 0 _0056_
rlabel metal2 40992 36232 40992 36232 0 _0057_
rlabel metal3 39592 36232 39592 36232 0 _0058_
rlabel metal2 39144 32312 39144 32312 0 _0059_
rlabel metal2 41496 33712 41496 33712 0 _0060_
rlabel metal2 35784 41048 35784 41048 0 _0061_
rlabel metal2 30968 35056 30968 35056 0 _0062_
rlabel metal3 19824 24920 19824 24920 0 _0063_
rlabel metal2 3304 45052 3304 45052 0 _0064_
rlabel metal2 7896 43064 7896 43064 0 _0065_
rlabel metal2 10360 46816 10360 46816 0 _0066_
rlabel metal2 7000 45864 7000 45864 0 _0067_
rlabel metal2 10920 45808 10920 45808 0 _0068_
rlabel metal2 9576 40992 9576 40992 0 _0069_
rlabel metal2 7672 48104 7672 48104 0 _0070_
rlabel metal3 10752 44296 10752 44296 0 _0071_
rlabel metal2 13832 41832 13832 41832 0 _0072_
rlabel metal2 12264 47432 12264 47432 0 _0073_
rlabel metal2 15624 42056 15624 42056 0 _0074_
rlabel metal3 25480 37352 25480 37352 0 _0075_
rlabel metal2 7000 45304 7000 45304 0 _0076_
rlabel metal2 7000 47600 7000 47600 0 _0077_
rlabel metal2 5376 41944 5376 41944 0 _0078_
rlabel metal3 6944 45752 6944 45752 0 _0079_
rlabel metal2 18088 42392 18088 42392 0 _0080_
rlabel metal2 15064 39816 15064 39816 0 _0081_
rlabel metal2 4200 45304 4200 45304 0 _0082_
rlabel metal2 6496 44520 6496 44520 0 _0083_
rlabel metal2 7112 37184 7112 37184 0 _0084_
rlabel metal2 14784 26488 14784 26488 0 _0085_
rlabel metal3 39032 35112 39032 35112 0 _0086_
rlabel metal2 12824 26824 12824 26824 0 _0087_
rlabel metal3 13720 25256 13720 25256 0 _0088_
rlabel metal2 18984 39424 18984 39424 0 _0089_
rlabel metal2 31528 39116 31528 39116 0 _0090_
rlabel metal2 34944 30184 34944 30184 0 _0091_
rlabel metal2 34328 30968 34328 30968 0 _0092_
rlabel metal2 32760 35672 32760 35672 0 _0093_
rlabel metal2 31808 39592 31808 39592 0 _0094_
rlabel metal2 4872 43568 4872 43568 0 _0095_
rlabel metal2 11928 40600 11928 40600 0 _0096_
rlabel metal2 12264 40768 12264 40768 0 _0097_
rlabel metal2 8232 39648 8232 39648 0 _0098_
rlabel metal2 7784 47096 7784 47096 0 _0099_
rlabel metal2 6776 40712 6776 40712 0 _0100_
rlabel metal2 2856 39872 2856 39872 0 _0101_
rlabel metal3 33320 39480 33320 39480 0 _0102_
rlabel metal2 32424 38780 32424 38780 0 _0103_
rlabel metal2 30800 38920 30800 38920 0 _0104_
rlabel metal2 17416 39648 17416 39648 0 _0105_
rlabel metal3 21504 42728 21504 42728 0 _0106_
rlabel metal2 15736 44128 15736 44128 0 _0107_
rlabel metal2 38472 30576 38472 30576 0 _0108_
rlabel metal2 38696 32872 38696 32872 0 _0109_
rlabel metal2 39480 31752 39480 31752 0 _0110_
rlabel metal3 33208 28056 33208 28056 0 _0111_
rlabel metal3 12040 24920 12040 24920 0 _0112_
rlabel metal2 29176 29008 29176 29008 0 _0113_
rlabel metal2 21784 42224 21784 42224 0 _0114_
rlabel metal3 26040 24920 26040 24920 0 _0115_
rlabel metal3 22176 24584 22176 24584 0 _0116_
rlabel metal3 34104 31528 34104 31528 0 _0117_
rlabel metal2 22568 36288 22568 36288 0 _0118_
rlabel metal2 9688 41888 9688 41888 0 _0119_
rlabel metal2 7952 39816 7952 39816 0 _0120_
rlabel metal2 19096 25704 19096 25704 0 _0121_
rlabel metal2 29288 28504 29288 28504 0 _0122_
rlabel metal2 30744 34496 30744 34496 0 _0123_
rlabel metal3 29008 29624 29008 29624 0 _0124_
rlabel metal2 27832 23968 27832 23968 0 _0125_
rlabel metal2 28280 26096 28280 26096 0 _0126_
rlabel metal2 11704 24360 11704 24360 0 _0127_
rlabel metal2 29624 29064 29624 29064 0 _0128_
rlabel metal2 21336 40320 21336 40320 0 _0129_
rlabel metal2 22008 32872 22008 32872 0 _0130_
rlabel metal3 10808 45080 10808 45080 0 _0131_
rlabel metal2 26152 31248 26152 31248 0 _0132_
rlabel metal2 26264 34160 26264 34160 0 _0133_
rlabel metal3 29064 29400 29064 29400 0 _0134_
rlabel metal2 25368 41776 25368 41776 0 _0135_
rlabel metal3 17304 32536 17304 32536 0 _0136_
rlabel metal3 21280 30072 21280 30072 0 _0137_
rlabel metal2 25144 30912 25144 30912 0 _0138_
rlabel metal2 25592 25816 25592 25816 0 _0139_
rlabel metal2 9688 34216 9688 34216 0 _0140_
rlabel metal2 22120 32648 22120 32648 0 _0141_
rlabel metal2 23520 37240 23520 37240 0 _0142_
rlabel metal2 25368 31696 25368 31696 0 _0143_
rlabel metal2 26824 32032 26824 32032 0 _0144_
rlabel metal3 19712 36344 19712 36344 0 _0145_
rlabel metal2 20104 28952 20104 28952 0 _0146_
rlabel metal2 8008 27720 8008 27720 0 _0147_
rlabel metal3 22176 30184 22176 30184 0 _0148_
rlabel metal2 24472 29344 24472 29344 0 _0149_
rlabel metal3 23072 29624 23072 29624 0 _0150_
rlabel metal2 27384 42336 27384 42336 0 _0151_
rlabel metal3 22120 42616 22120 42616 0 _0152_
rlabel metal2 13384 24752 13384 24752 0 _0153_
rlabel metal2 7896 25312 7896 25312 0 _0154_
rlabel metal2 13496 27832 13496 27832 0 _0155_
rlabel metal3 9408 43624 9408 43624 0 _0156_
rlabel metal2 8568 42392 8568 42392 0 _0157_
rlabel metal2 10248 49336 10248 49336 0 _0158_
rlabel metal3 14448 47432 14448 47432 0 _0159_
rlabel metal3 12320 43400 12320 43400 0 _0160_
rlabel metal2 16184 40600 16184 40600 0 _0161_
rlabel metal2 21672 47936 21672 47936 0 _0162_
rlabel metal2 15960 44632 15960 44632 0 _0163_
rlabel metal2 5992 42588 5992 42588 0 _0164_
rlabel metal3 6384 36344 6384 36344 0 _0165_
rlabel metal3 22680 31752 22680 31752 0 _0166_
rlabel metal2 20328 34048 20328 34048 0 _0167_
rlabel metal2 19544 39144 19544 39144 0 _0168_
rlabel metal2 16408 40880 16408 40880 0 _0169_
rlabel metal2 13608 46704 13608 46704 0 _0170_
rlabel metal2 14504 48216 14504 48216 0 _0171_
rlabel metal2 24472 24360 24472 24360 0 _0172_
rlabel metal3 6664 30128 6664 30128 0 _0173_
rlabel metal2 3864 45136 3864 45136 0 _0174_
rlabel metal3 7112 25704 7112 25704 0 _0175_
rlabel metal2 10808 39200 10808 39200 0 _0176_
rlabel metal3 20216 39144 20216 39144 0 _0177_
rlabel metal3 3080 39368 3080 39368 0 _0178_
rlabel metal2 3640 38528 3640 38528 0 _0179_
rlabel metal2 6440 29904 6440 29904 0 _0180_
rlabel metal2 6664 31304 6664 31304 0 _0181_
rlabel metal2 9016 29848 9016 29848 0 _0182_
rlabel metal2 21448 30800 21448 30800 0 _0183_
rlabel metal2 6888 40964 6888 40964 0 _0184_
rlabel metal2 7784 25144 7784 25144 0 _0185_
rlabel metal2 11312 26264 11312 26264 0 _0186_
rlabel metal2 11592 30352 11592 30352 0 _0187_
rlabel metal3 14224 34776 14224 34776 0 _0188_
rlabel metal2 19432 45528 19432 45528 0 _0189_
rlabel metal3 17192 42728 17192 42728 0 _0190_
rlabel metal1 24472 38696 24472 38696 0 _0191_
rlabel metal2 21672 44464 21672 44464 0 _0192_
rlabel metal2 18424 24416 18424 24416 0 _0193_
rlabel metal3 19320 44184 19320 44184 0 _0194_
rlabel metal3 17192 44184 17192 44184 0 _0195_
rlabel metal2 14728 24080 14728 24080 0 _0196_
rlabel metal2 23352 24920 23352 24920 0 _0197_
rlabel metal2 15904 27272 15904 27272 0 _0198_
rlabel metal2 14728 34440 14728 34440 0 _0199_
rlabel metal2 17192 27216 17192 27216 0 _0200_
rlabel metal2 15960 33712 15960 33712 0 _0201_
rlabel metal2 15848 34552 15848 34552 0 _0202_
rlabel metal2 17192 39900 17192 39900 0 _0203_
rlabel metal2 3248 31752 3248 31752 0 _0204_
rlabel metal2 2968 30240 2968 30240 0 _0205_
rlabel metal2 5320 40264 5320 40264 0 _0206_
rlabel metal2 3304 30296 3304 30296 0 _0207_
rlabel metal2 34104 39592 34104 39592 0 _0208_
rlabel metal3 31192 40376 31192 40376 0 _0209_
rlabel metal3 13832 46648 13832 46648 0 _0210_
rlabel metal2 31416 39816 31416 39816 0 _0211_
rlabel metal2 5824 23240 5824 23240 0 _0212_
rlabel metal2 7448 32256 7448 32256 0 _0213_
rlabel metal2 12040 35560 12040 35560 0 _0214_
rlabel metal3 17920 30968 17920 30968 0 _0215_
rlabel metal2 4872 31640 4872 31640 0 _0216_
rlabel metal2 2632 39200 2632 39200 0 _0217_
rlabel metal2 2464 38024 2464 38024 0 _0218_
rlabel metal2 3080 34552 3080 34552 0 _0219_
rlabel metal3 5544 33320 5544 33320 0 _0220_
rlabel metal2 15400 27720 15400 27720 0 _0221_
rlabel metal3 12040 43512 12040 43512 0 _0222_
rlabel metal2 21560 37408 21560 37408 0 _0223_
rlabel metal2 24696 27664 24696 27664 0 _0224_
rlabel metal2 23632 42840 23632 42840 0 _0225_
rlabel metal2 14056 24584 14056 24584 0 _0226_
rlabel metal2 8680 29400 8680 29400 0 _0227_
rlabel metal2 8792 28224 8792 28224 0 _0228_
rlabel metal3 15876 31752 15876 31752 0 _0229_
rlabel metal2 15736 40936 15736 40936 0 _0230_
rlabel metal3 26880 47488 26880 47488 0 _0231_
rlabel metal2 18648 25144 18648 25144 0 _0232_
rlabel metal2 19208 22904 19208 22904 0 _0233_
rlabel metal3 17304 24696 17304 24696 0 _0234_
rlabel metal2 22120 23912 22120 23912 0 _0235_
rlabel metal2 18648 44744 18648 44744 0 _0236_
rlabel metal2 9912 24640 9912 24640 0 _0237_
rlabel metal2 21112 24248 21112 24248 0 _0238_
rlabel metal2 14504 44968 14504 44968 0 _0239_
rlabel metal2 20440 25088 20440 25088 0 _0240_
rlabel metal2 23688 42224 23688 42224 0 _0241_
rlabel metal3 17808 33208 17808 33208 0 _0242_
rlabel metal2 22680 25760 22680 25760 0 _0243_
rlabel metal2 18032 36344 18032 36344 0 _0244_
rlabel metal2 20832 33096 20832 33096 0 _0245_
rlabel metal2 23016 35616 23016 35616 0 _0246_
rlabel metal3 8148 26376 8148 26376 0 _0247_
rlabel metal2 23464 26236 23464 26236 0 _0248_
rlabel metal2 7728 37240 7728 37240 0 _0249_
rlabel metal2 8568 34664 8568 34664 0 _0250_
rlabel metal2 25816 36736 25816 36736 0 _0251_
rlabel metal2 23912 36008 23912 36008 0 _0252_
rlabel metal2 23464 36232 23464 36232 0 _0253_
rlabel metal3 18816 36232 18816 36232 0 _0254_
rlabel metal2 20328 35168 20328 35168 0 _0255_
rlabel metal2 21000 34272 21000 34272 0 _0256_
rlabel metal2 21560 34944 21560 34944 0 _0257_
rlabel metal2 18984 37912 18984 37912 0 _0258_
rlabel metal2 13160 31248 13160 31248 0 _0259_
rlabel metal2 15176 31472 15176 31472 0 _0260_
rlabel metal2 18536 34608 18536 34608 0 _0261_
rlabel metal2 25256 36400 25256 36400 0 _0262_
rlabel metal3 25200 39256 25200 39256 0 _0263_
rlabel metal2 27160 47628 27160 47628 0 _0264_
rlabel metal2 11816 39648 11816 39648 0 _0265_
rlabel metal2 16016 28616 16016 28616 0 _0266_
rlabel metal3 22624 27832 22624 27832 0 _0267_
rlabel metal2 24696 44800 24696 44800 0 _0268_
rlabel metal2 25480 37296 25480 37296 0 _0269_
rlabel metal4 26152 40040 26152 40040 0 _0270_
rlabel metal3 8904 25480 8904 25480 0 _0271_
rlabel metal2 9184 32760 9184 32760 0 _0272_
rlabel metal2 10472 25424 10472 25424 0 _0273_
rlabel metal3 11704 25368 11704 25368 0 _0274_
rlabel metal2 12040 26040 12040 26040 0 _0275_
rlabel metal2 12040 47768 12040 47768 0 _0276_
rlabel metal2 11816 26152 11816 26152 0 _0277_
rlabel metal3 11480 25480 11480 25480 0 _0278_
rlabel metal2 11368 24696 11368 24696 0 _0279_
rlabel metal2 24472 45080 24472 45080 0 _0280_
rlabel metal2 27160 45024 27160 45024 0 _0281_
rlabel metal3 27832 48216 27832 48216 0 _0282_
rlabel metal3 27328 45192 27328 45192 0 _0283_
rlabel metal2 30072 45080 30072 45080 0 _0284_
rlabel metal2 16184 50344 16184 50344 0 _0285_
rlabel metal2 15512 48104 15512 48104 0 _0286_
rlabel metal2 23240 41216 23240 41216 0 _0287_
rlabel metal3 18648 33992 18648 33992 0 _0288_
rlabel metal2 16184 45024 16184 45024 0 _0289_
rlabel metal2 18200 47600 18200 47600 0 _0290_
rlabel metal2 17192 47712 17192 47712 0 _0291_
rlabel metal2 17416 43792 17416 43792 0 _0292_
rlabel metal2 18536 32256 18536 32256 0 _0293_
rlabel metal2 17360 41384 17360 41384 0 _0294_
rlabel metal2 17528 40544 17528 40544 0 _0295_
rlabel metal2 16408 44016 16408 44016 0 _0296_
rlabel metal2 2632 33096 2632 33096 0 _0297_
rlabel metal3 4480 35672 4480 35672 0 _0298_
rlabel metal2 3920 33320 3920 33320 0 _0299_
rlabel metal3 15876 44296 15876 44296 0 _0300_
rlabel metal2 18144 30968 18144 30968 0 _0301_
rlabel metal3 13048 34888 13048 34888 0 _0302_
rlabel metal2 15176 31808 15176 31808 0 _0303_
rlabel metal2 16296 30856 16296 30856 0 _0304_
rlabel metal2 19096 32144 19096 32144 0 _0305_
rlabel metal2 16688 39368 16688 39368 0 _0306_
rlabel metal3 17472 44296 17472 44296 0 _0307_
rlabel metal3 17528 44072 17528 44072 0 _0308_
rlabel metal2 30072 37184 30072 37184 0 _0309_
rlabel metal2 29792 37464 29792 37464 0 _0310_
rlabel metal2 28728 37184 28728 37184 0 _0311_
rlabel metal3 26992 38696 26992 38696 0 _0312_
rlabel metal2 13048 41216 13048 41216 0 _0313_
rlabel metal2 26152 40152 26152 40152 0 _0314_
rlabel metal2 25200 33208 25200 33208 0 _0315_
rlabel metal2 22792 25312 22792 25312 0 _0316_
rlabel metal2 25816 39088 25816 39088 0 _0317_
rlabel metal2 12376 36456 12376 36456 0 _0318_
rlabel metal3 19992 37352 19992 37352 0 _0319_
rlabel metal3 19992 38080 19992 38080 0 _0320_
rlabel metal3 18032 41048 18032 41048 0 _0321_
rlabel metal3 24640 38696 24640 38696 0 _0322_
rlabel metal3 25536 39032 25536 39032 0 _0323_
rlabel metal2 27496 48328 27496 48328 0 _0324_
rlabel metal3 25144 49000 25144 49000 0 _0325_
rlabel metal3 24304 33432 24304 33432 0 _0326_
rlabel metal3 25984 39256 25984 39256 0 _0327_
rlabel metal2 27720 35448 27720 35448 0 _0328_
rlabel metal2 28056 34272 28056 34272 0 _0329_
rlabel metal2 28504 40376 28504 40376 0 _0330_
rlabel metal2 27944 40040 27944 40040 0 _0331_
rlabel metal2 2912 34776 2912 34776 0 _0332_
rlabel metal2 18760 40544 18760 40544 0 _0333_
rlabel metal2 18648 38668 18648 38668 0 _0334_
rlabel metal2 18704 37464 18704 37464 0 _0335_
rlabel metal2 19096 37072 19096 37072 0 _0336_
rlabel metal2 19320 34552 19320 34552 0 _0337_
rlabel metal2 17304 37632 17304 37632 0 _0338_
rlabel metal2 17640 34048 17640 34048 0 _0339_
rlabel metal2 17304 38024 17304 38024 0 _0340_
rlabel metal3 18200 38024 18200 38024 0 _0341_
rlabel metal2 19208 30296 19208 30296 0 _0342_
rlabel metal2 18760 28728 18760 28728 0 _0343_
rlabel metal2 18256 28056 18256 28056 0 _0344_
rlabel metal3 18592 23240 18592 23240 0 _0345_
rlabel metal2 18872 27832 18872 27832 0 _0346_
rlabel metal2 18424 27272 18424 27272 0 _0347_
rlabel metal3 10640 26376 10640 26376 0 _0348_
rlabel metal2 9856 26488 9856 26488 0 _0349_
rlabel metal2 17752 27160 17752 27160 0 _0350_
rlabel metal2 18256 32088 18256 32088 0 _0351_
rlabel metal2 18984 38248 18984 38248 0 _0352_
rlabel metal2 17864 42224 17864 42224 0 _0353_
rlabel metal3 19208 41944 19208 41944 0 _0354_
rlabel metal2 19656 41440 19656 41440 0 _0355_
rlabel metal2 18480 47656 18480 47656 0 _0356_
rlabel metal2 18592 41944 18592 41944 0 _0357_
rlabel metal2 18704 39368 18704 39368 0 _0358_
rlabel metal2 19096 41048 19096 41048 0 _0359_
rlabel metal2 19544 40880 19544 40880 0 _0360_
rlabel metal3 25984 45752 25984 45752 0 _0361_
rlabel metal3 28504 37128 28504 37128 0 _0362_
rlabel metal2 27440 37016 27440 37016 0 _0363_
rlabel metal2 27832 31808 27832 31808 0 _0364_
rlabel metal2 17976 31024 17976 31024 0 _0365_
rlabel metal2 28056 31192 28056 31192 0 _0366_
rlabel metal2 27832 43512 27832 43512 0 _0367_
rlabel metal4 26824 41664 26824 41664 0 _0368_
rlabel metal2 5432 26264 5432 26264 0 _0369_
rlabel metal2 8904 33376 8904 33376 0 _0370_
rlabel metal3 15960 26488 15960 26488 0 _0371_
rlabel metal2 22512 40936 22512 40936 0 _0372_
rlabel metal2 14392 29344 14392 29344 0 _0373_
rlabel metal2 15064 28840 15064 28840 0 _0374_
rlabel metal2 14728 29624 14728 29624 0 _0375_
rlabel metal3 20160 40376 20160 40376 0 _0376_
rlabel metal2 24808 44464 24808 44464 0 _0377_
rlabel metal2 22456 48048 22456 48048 0 _0378_
rlabel metal2 22792 47936 22792 47936 0 _0379_
rlabel metal2 23912 48384 23912 48384 0 _0380_
rlabel metal2 24024 47432 24024 47432 0 _0381_
rlabel metal2 27832 47432 27832 47432 0 _0382_
rlabel metal2 27720 48496 27720 48496 0 _0383_
rlabel metal3 24696 43232 24696 43232 0 _0384_
rlabel metal2 24024 43288 24024 43288 0 _0385_
rlabel metal2 28280 44912 28280 44912 0 _0386_
rlabel metal2 25032 43176 25032 43176 0 _0387_
rlabel metal3 25032 28056 25032 28056 0 _0388_
rlabel metal3 21672 31080 21672 31080 0 _0389_
rlabel metal3 25256 30968 25256 30968 0 _0390_
rlabel metal3 26040 40152 26040 40152 0 _0391_
rlabel metal2 25256 41272 25256 41272 0 _0392_
rlabel metal3 20216 23408 20216 23408 0 _0393_
rlabel metal2 10360 31752 10360 31752 0 _0394_
rlabel metal3 9240 28056 9240 28056 0 _0395_
rlabel metal2 10752 28728 10752 28728 0 _0396_
rlabel metal2 10248 28896 10248 28896 0 _0397_
rlabel metal2 5656 30296 5656 30296 0 _0398_
rlabel metal3 3920 30856 3920 30856 0 _0399_
rlabel metal2 6328 29736 6328 29736 0 _0400_
rlabel metal2 2520 41496 2520 41496 0 _0401_
rlabel metal3 2352 44856 2352 44856 0 _0402_
rlabel metal2 14728 25424 14728 25424 0 _0403_
rlabel metal3 14224 26824 14224 26824 0 _0404_
rlabel metal3 8008 27160 8008 27160 0 _0405_
rlabel metal3 7896 26488 7896 26488 0 _0406_
rlabel metal2 5432 27776 5432 27776 0 _0407_
rlabel metal2 7168 28056 7168 28056 0 _0408_
rlabel metal2 8008 24192 8008 24192 0 _0409_
rlabel metal3 20888 34664 20888 34664 0 _0410_
rlabel metal2 21224 38724 21224 38724 0 _0411_
rlabel metal2 23464 42616 23464 42616 0 _0412_
rlabel metal2 18536 49784 18536 49784 0 _0413_
rlabel metal2 19096 49056 19096 49056 0 _0414_
rlabel metal2 25816 43904 25816 43904 0 _0415_
rlabel metal2 26264 43792 26264 43792 0 _0416_
rlabel metal3 35224 45864 35224 45864 0 _0417_
rlabel metal2 32984 41888 32984 41888 0 _0418_
rlabel metal2 19656 47432 19656 47432 0 _0419_
rlabel metal2 22064 44856 22064 44856 0 _0420_
rlabel metal2 22904 45192 22904 45192 0 _0421_
rlabel metal2 19320 28840 19320 28840 0 _0422_
rlabel metal2 18760 35336 18760 35336 0 _0423_
rlabel metal2 15736 26656 15736 26656 0 _0424_
rlabel metal4 17640 33152 17640 33152 0 _0425_
rlabel metal3 3920 32088 3920 32088 0 _0426_
rlabel metal2 3472 35896 3472 35896 0 _0427_
rlabel metal2 2912 35000 2912 35000 0 _0428_
rlabel metal3 17752 35896 17752 35896 0 _0429_
rlabel metal2 23128 44464 23128 44464 0 _0430_
rlabel metal2 29400 45584 29400 45584 0 _0431_
rlabel metal2 26488 33544 26488 33544 0 _0432_
rlabel metal2 29960 39368 29960 39368 0 _0433_
rlabel metal2 26768 40600 26768 40600 0 _0434_
rlabel metal2 29512 43960 29512 43960 0 _0435_
rlabel metal2 40936 41440 40936 41440 0 _0436_
rlabel metal2 26600 38472 26600 38472 0 _0437_
rlabel metal2 23464 41048 23464 41048 0 _0438_
rlabel metal2 21336 39144 21336 39144 0 _0439_
rlabel metal2 20384 36456 20384 36456 0 _0440_
rlabel metal2 20776 38808 20776 38808 0 _0441_
rlabel metal3 24472 38808 24472 38808 0 _0442_
rlabel metal3 13160 39144 13160 39144 0 _0443_
rlabel metal3 8904 29960 8904 29960 0 _0444_
rlabel metal2 3640 36904 3640 36904 0 _0445_
rlabel metal3 18872 38752 18872 38752 0 _0446_
rlabel metal2 27608 39088 27608 39088 0 _0447_
rlabel metal2 20832 24136 20832 24136 0 _0448_
rlabel metal2 15288 26908 15288 26908 0 _0449_
rlabel metal2 15848 27720 15848 27720 0 _0450_
rlabel metal2 19656 48552 19656 48552 0 _0451_
rlabel metal2 27048 39480 27048 39480 0 _0452_
rlabel metal2 18088 24752 18088 24752 0 _0453_
rlabel metal2 16184 23408 16184 23408 0 _0454_
rlabel metal2 16576 25592 16576 25592 0 _0455_
rlabel metal3 20160 24024 20160 24024 0 _0456_
rlabel metal2 23240 48216 23240 48216 0 _0457_
rlabel metal4 23688 42784 23688 42784 0 _0458_
rlabel metal2 26488 40376 26488 40376 0 _0459_
rlabel metal3 36064 42728 36064 42728 0 _0460_
rlabel metal3 28840 42728 28840 42728 0 _0461_
rlabel metal2 29960 43792 29960 43792 0 _0462_
rlabel metal3 21336 41384 21336 41384 0 _0463_
rlabel metal2 21504 39592 21504 39592 0 _0464_
rlabel metal2 21560 30632 21560 30632 0 _0465_
rlabel metal3 20720 29624 20720 29624 0 _0466_
rlabel metal3 21616 41160 21616 41160 0 _0467_
rlabel metal2 22120 41664 22120 41664 0 _0468_
rlabel metal3 13216 38360 13216 38360 0 _0469_
rlabel metal2 4088 39536 4088 39536 0 _0470_
rlabel metal2 4200 36456 4200 36456 0 _0471_
rlabel metal2 8232 37744 8232 37744 0 _0472_
rlabel metal2 22232 41888 22232 41888 0 _0473_
rlabel metal2 21560 45864 21560 45864 0 _0474_
rlabel metal2 21504 45304 21504 45304 0 _0475_
rlabel metal2 22456 43792 22456 43792 0 _0476_
rlabel metal2 22904 42056 22904 42056 0 _0477_
rlabel metal2 33320 44240 33320 44240 0 _0478_
rlabel metal2 30072 42056 30072 42056 0 _0479_
rlabel metal2 30072 43624 30072 43624 0 _0480_
rlabel metal2 19320 47992 19320 47992 0 _0481_
rlabel metal2 20104 48328 20104 48328 0 _0482_
rlabel metal2 20328 47768 20328 47768 0 _0483_
rlabel metal2 12936 30576 12936 30576 0 _0484_
rlabel metal3 14560 36680 14560 36680 0 _0485_
rlabel metal2 16072 36568 16072 36568 0 _0486_
rlabel metal2 15176 37296 15176 37296 0 _0487_
rlabel metal2 15456 38584 15456 38584 0 _0488_
rlabel metal2 16576 39256 16576 39256 0 _0489_
rlabel metal2 2856 43008 2856 43008 0 _0490_
rlabel metal2 3136 40600 3136 40600 0 _0491_
rlabel metal2 18760 43288 18760 43288 0 _0492_
rlabel metal2 30632 43960 30632 43960 0 _0493_
rlabel metal3 29456 54488 29456 54488 0 _0494_
rlabel metal3 10248 53032 10248 53032 0 _0495_
rlabel metal2 12488 54880 12488 54880 0 _0496_
rlabel metal2 12376 53088 12376 53088 0 _0497_
rlabel via2 11704 52696 11704 52696 0 _0498_
rlabel metal2 12600 50176 12600 50176 0 _0499_
rlabel metal2 11256 50876 11256 50876 0 _0500_
rlabel metal2 29288 53312 29288 53312 0 _0501_
rlabel metal3 11200 51464 11200 51464 0 _0502_
rlabel metal2 27608 54712 27608 54712 0 _0503_
rlabel metal2 11424 50456 11424 50456 0 _0504_
rlabel metal2 29624 52360 29624 52360 0 _0505_
rlabel metal2 13776 44408 13776 44408 0 _0506_
rlabel metal2 11928 52248 11928 52248 0 _0507_
rlabel metal2 32592 53816 32592 53816 0 _0508_
rlabel metal2 35000 43904 35000 43904 0 _0509_
rlabel metal2 34440 45640 34440 45640 0 _0510_
rlabel metal2 36008 41608 36008 41608 0 _0511_
rlabel metal3 37744 53144 37744 53144 0 _0512_
rlabel metal2 34664 40432 34664 40432 0 _0513_
rlabel metal3 39312 51464 39312 51464 0 _0514_
rlabel metal2 35784 41440 35784 41440 0 _0515_
rlabel metal3 40880 54712 40880 54712 0 _0516_
rlabel metal3 33880 44296 33880 44296 0 _0517_
rlabel metal2 38920 47152 38920 47152 0 _0518_
rlabel metal2 22456 50624 22456 50624 0 _0519_
rlabel metal2 24696 50456 24696 50456 0 _0520_
rlabel metal3 28000 52808 28000 52808 0 _0521_
rlabel metal2 24024 51968 24024 51968 0 _0522_
rlabel metal3 23352 50680 23352 50680 0 _0523_
rlabel metal3 25816 53592 25816 53592 0 _0524_
rlabel metal3 23296 53816 23296 53816 0 _0525_
rlabel metal3 26432 50568 26432 50568 0 _0526_
rlabel metal2 41944 46312 41944 46312 0 _0527_
rlabel metal2 39480 45920 39480 45920 0 _0528_
rlabel metal2 39480 47096 39480 47096 0 _0529_
rlabel metal2 40936 46816 40936 46816 0 _0530_
rlabel metal2 40824 43204 40824 43204 0 _0531_
rlabel metal2 39088 42840 39088 42840 0 _0532_
rlabel metal2 40264 45528 40264 45528 0 _0533_
rlabel metal2 29848 53760 29848 53760 0 _0534_
rlabel metal2 30408 54040 30408 54040 0 _0535_
rlabel metal2 36400 54712 36400 54712 0 _0536_
rlabel metal2 31752 54432 31752 54432 0 _0537_
rlabel metal2 30856 52864 30856 52864 0 _0538_
rlabel metal2 33992 54432 33992 54432 0 _0539_
rlabel metal2 42336 53480 42336 53480 0 _0540_
rlabel metal3 35896 52920 35896 52920 0 _0541_
rlabel metal3 40320 54600 40320 54600 0 _0542_
rlabel metal2 41720 53312 41720 53312 0 _0543_
rlabel metal2 39592 51296 39592 51296 0 _0544_
rlabel metal2 41944 52416 41944 52416 0 _0545_
rlabel metal2 41832 51296 41832 51296 0 _0546_
rlabel metal2 41048 54152 41048 54152 0 _0547_
rlabel metal2 30408 50848 30408 50848 0 _0548_
rlabel metal2 14616 53312 14616 53312 0 _0549_
rlabel metal2 15624 52192 15624 52192 0 _0550_
rlabel metal3 17472 52136 17472 52136 0 _0551_
rlabel metal2 15288 54656 15288 54656 0 _0552_
rlabel metal3 15456 51912 15456 51912 0 _0553_
rlabel metal3 18144 54488 18144 54488 0 _0554_
rlabel metal2 18312 51856 18312 51856 0 _0555_
rlabel metal2 35224 47432 35224 47432 0 _0556_
rlabel metal3 31920 50008 31920 50008 0 _0557_
rlabel metal2 33768 48608 33768 48608 0 _0558_
rlabel metal2 32872 46312 32872 46312 0 _0559_
rlabel metal2 34384 47544 34384 47544 0 _0560_
rlabel metal2 34776 46648 34776 46648 0 _0561_
rlabel metal2 31808 48328 31808 48328 0 _0562_
rlabel metal2 23128 57778 23128 57778 0 bus_in[0]
rlabel metal2 25368 57778 25368 57778 0 bus_in[1]
rlabel metal2 27944 56728 27944 56728 0 bus_in[2]
rlabel metal2 29848 57778 29848 57778 0 bus_in[3]
rlabel metal2 32088 57778 32088 57778 0 bus_in[4]
rlabel metal2 34328 57778 34328 57778 0 bus_in[5]
rlabel metal2 36568 57778 36568 57778 0 bus_in[6]
rlabel metal2 39368 56448 39368 56448 0 bus_in[7]
rlabel metal2 41048 57778 41048 57778 0 bus_out[0]
rlabel metal2 43288 57778 43288 57778 0 bus_out[1]
rlabel metal3 46144 55384 46144 55384 0 bus_out[2]
rlabel metal2 47768 57778 47768 57778 0 bus_out[3]
rlabel metal2 50008 57778 50008 57778 0 bus_out[4]
rlabel metal3 53032 55384 53032 55384 0 bus_out[5]
rlabel metal2 54488 57778 54488 57778 0 bus_out[6]
rlabel metal2 56728 57330 56728 57330 0 bus_out[7]
rlabel metal2 27496 52136 27496 52136 0 clknet_0_wb_clk_i
rlabel metal2 25256 52080 25256 52080 0 clknet_2_0__leaf_wb_clk_i
rlabel metal3 6048 51352 6048 51352 0 clknet_2_1__leaf_wb_clk_i
rlabel metal2 41104 42728 41104 42728 0 clknet_2_2__leaf_wb_clk_i
rlabel metal3 33432 55272 33432 55272 0 clknet_2_3__leaf_wb_clk_i
rlabel metal2 16464 56280 16464 56280 0 cs_port[0]
rlabel metal2 18648 57778 18648 57778 0 cs_port[1]
rlabel metal2 21000 56168 21000 56168 0 cs_port[2]
rlabel metal2 2184 48552 2184 48552 0 full_addr\[0\]
rlabel metal2 36680 54992 36680 54992 0 full_addr\[10\]
rlabel metal2 36568 52864 36568 52864 0 full_addr\[11\]
rlabel metal2 40264 51800 40264 51800 0 full_addr\[12\]
rlabel metal2 42728 52416 42728 52416 0 full_addr\[13\]
rlabel metal2 42504 50904 42504 50904 0 full_addr\[14\]
rlabel metal2 43120 52136 43120 52136 0 full_addr\[15\]
rlabel metal3 2520 50680 2520 50680 0 full_addr\[1\]
rlabel metal3 6608 50792 6608 50792 0 full_addr\[2\]
rlabel metal2 7112 50960 7112 50960 0 full_addr\[3\]
rlabel metal2 39928 39256 39928 39256 0 full_addr\[4\]
rlabel metal2 38696 36848 38696 36848 0 full_addr\[5\]
rlabel metal2 40264 38024 40264 38024 0 full_addr\[6\]
rlabel metal2 40376 35952 40376 35952 0 full_addr\[7\]
rlabel metal2 32088 53984 32088 53984 0 full_addr\[8\]
rlabel metal3 34552 53032 34552 53032 0 full_addr\[9\]
rlabel metal2 11928 57778 11928 57778 0 le_hi_act
rlabel metal2 9688 57778 9688 57778 0 le_lo_act
rlabel metal2 8120 55440 8120 55440 0 net1
rlabel metal2 18200 47992 18200 47992 0 net10
rlabel metal2 18648 48160 18648 48160 0 net11
rlabel metal2 20104 46256 20104 46256 0 net12
rlabel metal2 29176 54656 29176 54656 0 net13
rlabel metal2 10248 52752 10248 52752 0 net14
rlabel metal3 4144 30072 4144 30072 0 net15
rlabel metal2 1848 42280 1848 42280 0 net16
rlabel metal3 2408 51464 2408 51464 0 net17
rlabel metal2 2184 53032 2184 53032 0 net18
rlabel metal3 1736 54600 1736 54600 0 net19
rlabel metal2 23016 55440 23016 55440 0 net2
rlabel metal2 2016 55440 2016 55440 0 net20
rlabel metal2 2520 55440 2520 55440 0 net21
rlabel metal3 2856 33096 2856 33096 0 net22
rlabel metal2 6552 33376 6552 33376 0 net23
rlabel metal2 2072 37016 2072 37016 0 net24
rlabel metal2 2744 34832 2744 34832 0 net25
rlabel metal3 1624 39592 1624 39592 0 net26
rlabel metal2 2072 41496 2072 41496 0 net27
rlabel metal2 2072 43008 2072 43008 0 net28
rlabel metal2 2408 39144 2408 39144 0 net29
rlabel metal2 25424 55272 25424 55272 0 net3
rlabel metal2 2072 42392 2072 42392 0 net30
rlabel metal2 2352 3640 2352 3640 0 net31
rlabel metal2 2072 21280 2072 21280 0 net32
rlabel metal2 2016 22232 2016 22232 0 net33
rlabel metal3 2632 23800 2632 23800 0 net34
rlabel metal2 2128 25368 2128 25368 0 net35
rlabel metal2 2072 28280 2072 28280 0 net36
rlabel metal2 2800 28616 2800 28616 0 net37
rlabel metal3 5152 4536 5152 4536 0 net38
rlabel metal2 2184 5824 2184 5824 0 net39
rlabel metal2 27720 55356 27720 55356 0 net4
rlabel metal2 4816 25032 4816 25032 0 net40
rlabel metal2 2016 9688 2016 9688 0 net41
rlabel metal3 4200 11256 4200 11256 0 net42
rlabel metal2 2072 13104 2072 13104 0 net43
rlabel metal2 1960 15512 1960 15512 0 net44
rlabel metal2 2072 22008 2072 22008 0 net45
rlabel metal3 1736 23464 1736 23464 0 net46
rlabel metal2 13720 54964 13720 54964 0 net47
rlabel metal2 5880 55664 5880 55664 0 net48
rlabel metal2 30576 53928 30576 53928 0 net49
rlabel metal2 29736 53592 29736 53592 0 net5
rlabel metal2 43736 55552 43736 55552 0 net50
rlabel metal2 45416 51968 45416 51968 0 net51
rlabel metal2 47880 56056 47880 56056 0 net52
rlabel metal2 50904 54432 50904 54432 0 net53
rlabel metal2 52696 55160 52696 55160 0 net54
rlabel metal3 49616 53816 49616 53816 0 net55
rlabel metal2 55384 49392 55384 49392 0 net56
rlabel metal2 32648 55720 32648 55720 0 net6
rlabel metal2 34832 54600 34832 54600 0 net7
rlabel metal2 37128 55720 37128 55720 0 net8
rlabel metal2 39256 55412 39256 55412 0 net9
rlabel metal2 1736 30464 1736 30464 0 ram_end[0]
rlabel metal2 1736 48776 1736 48776 0 ram_end[10]
rlabel metal2 1848 50904 1848 50904 0 ram_end[11]
rlabel metal2 1736 52584 1736 52584 0 ram_end[12]
rlabel metal2 1736 54264 1736 54264 0 ram_end[13]
rlabel metal2 1736 55944 1736 55944 0 ram_end[14]
rlabel metal3 1470 57624 1470 57624 0 ram_end[15]
rlabel metal2 1736 32872 1736 32872 0 ram_end[1]
rlabel metal3 1246 34328 1246 34328 0 ram_end[2]
rlabel metal2 1736 36680 1736 36680 0 ram_end[3]
rlabel metal2 1848 38668 1848 38668 0 ram_end[4]
rlabel metal2 1736 40040 1736 40040 0 ram_end[5]
rlabel metal2 1736 41328 1736 41328 0 ram_end[6]
rlabel metal2 1848 43344 1848 43344 0 ram_end[7]
rlabel metal2 1736 45416 1736 45416 0 ram_end[8]
rlabel metal2 1736 46816 1736 46816 0 ram_end[9]
rlabel metal2 1736 2744 1736 2744 0 ram_start[0]
rlabel metal3 1246 19992 1246 19992 0 ram_start[10]
rlabel metal2 1736 22008 1736 22008 0 ram_start[11]
rlabel metal2 1736 23688 1736 23688 0 ram_start[12]
rlabel metal3 1246 25368 1246 25368 0 ram_start[13]
rlabel metal2 1736 27496 1736 27496 0 ram_start[14]
rlabel metal2 2408 29512 2408 29512 0 ram_start[15]
rlabel metal2 1736 4088 1736 4088 0 ram_start[1]
rlabel metal2 1736 5768 1736 5768 0 ram_start[2]
rlabel metal2 1736 7784 1736 7784 0 ram_start[3]
rlabel metal2 1736 9464 1736 9464 0 ram_start[4]
rlabel metal2 1736 11144 1736 11144 0 ram_start[5]
rlabel metal3 1246 12824 1246 12824 0 ram_start[6]
rlabel metal2 1736 14952 1736 14952 0 ram_start[7]
rlabel metal2 1736 16632 1736 16632 0 ram_start[8]
rlabel metal2 1736 18312 1736 18312 0 ram_start[9]
rlabel metal2 14168 57778 14168 57778 0 rom_enabled
rlabel metal2 5152 56280 5152 56280 0 rst
rlabel metal3 4368 53816 4368 53816 0 wb_clk_i
rlabel metal3 24528 49896 24528 49896 0 writable\[0\]
rlabel metal2 23016 49224 23016 49224 0 writable\[10\]
rlabel metal3 20328 49896 20328 49896 0 writable\[11\]
rlabel metal3 22568 46928 22568 46928 0 writable\[12\]
rlabel metal2 22904 48552 22904 48552 0 writable\[13\]
rlabel metal2 22680 46088 22680 46088 0 writable\[14\]
rlabel metal3 23660 48888 23660 48888 0 writable\[15\]
rlabel metal2 28168 54096 28168 54096 0 writable\[1\]
rlabel metal2 24528 49112 24528 49112 0 writable\[2\]
rlabel metal2 25928 52080 25928 52080 0 writable\[3\]
rlabel metal2 39256 47096 39256 47096 0 writable\[4\]
rlabel metal2 41384 43176 41384 43176 0 writable\[5\]
rlabel metal2 38696 43120 38696 43120 0 writable\[6\]
rlabel metal2 40152 45024 40152 45024 0 writable\[7\]
rlabel metal2 15960 53872 15960 53872 0 writable\[8\]
rlabel metal2 16016 51240 16016 51240 0 writable\[9\]
<< properties >>
string FIXED_BBOX 0 0 60000 60000
<< end >>
